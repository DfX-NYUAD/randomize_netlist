// Randomized netlist
//
// Parameter ``netlist.v'': b14_original_6_metal_layers.v
// Parameter ``cells.inputs'': cells.inputs
// Parameter ``cells.outputs'': cells.outputs
// Parameter ``cells.functions'': cells.functions
// Parameter ``golden_netlist'': b14_original_6_metal_layers.v
// Parameter ``also_output_scrambled_netlists'': 0
// Parameter ``threads'': 32
// Parameter ``intermediate_output_HD_step'': 0.05
// Parameter ``HD_target'': 0.5
// Parameter ``acceptance_ratio'': 0.01
// Parameter ``HD_sampling_iterations'': 1,000
// Parameter ``lazy_Boolean_evaluation'': 0
// Parameter ``consider_fanout'': 0
// Parameter ``consider_driving_strength'': 1
// Parameter ``random_op'': -1
//  Replace underlying cell type: 1
//  Swap outputs for a pair of gates: 2
//  Swap inputs for a pair of gates: 3
//  Delete a gate: 4
//  Insert a gate: 5
//  Randomly any of the above operation: -1
//
//
// Achieved the following HD for this randomized netlist: 0.0585818
//
// Randomization iterations: 41
//
// Replaced cell type for that many gates: 3
// Swapped outputs for that many pairs of gates: 3
// Swapped inputs for that many pairs of gates: 2
// Deleted that many gates: 4
// Inserted that many gates: 8
//

module b14_rand (
DATAI_31_,
DATAI_30_,
DATAI_29_,
DATAI_28_,
DATAI_27_,
DATAI_26_,
DATAI_25_,
DATAI_24_,
DATAI_23_,
DATAI_22_,
DATAI_21_,
DATAI_20_,
DATAI_19_,
DATAI_18_,
DATAI_17_,
DATAI_16_,
DATAI_15_,
DATAI_14_,
DATAI_13_,
DATAI_12_,
DATAI_11_,
DATAI_10_,
DATAI_9_,
DATAI_8_,
DATAI_7_,
DATAI_6_,
DATAI_5_,
DATAI_4_,
DATAI_3_,
DATAI_2_,
DATAI_1_,
DATAI_0_,
STATE_REG_SCAN_IN,
REG3_REG_7__SCAN_IN,
REG3_REG_27__SCAN_IN,
REG3_REG_14__SCAN_IN,
REG3_REG_23__SCAN_IN,
REG3_REG_10__SCAN_IN,
REG3_REG_3__SCAN_IN,
REG3_REG_19__SCAN_IN,
REG3_REG_28__SCAN_IN,
REG3_REG_8__SCAN_IN,
REG3_REG_1__SCAN_IN,
REG3_REG_21__SCAN_IN,
REG3_REG_12__SCAN_IN,
REG3_REG_25__SCAN_IN,
REG3_REG_16__SCAN_IN,
REG3_REG_5__SCAN_IN,
REG3_REG_17__SCAN_IN,
REG3_REG_24__SCAN_IN,
REG3_REG_4__SCAN_IN,
REG3_REG_9__SCAN_IN,
REG3_REG_0__SCAN_IN,
REG3_REG_20__SCAN_IN,
REG3_REG_13__SCAN_IN,
IR_REG_0__SCAN_IN,
IR_REG_1__SCAN_IN,
IR_REG_2__SCAN_IN,
IR_REG_3__SCAN_IN,
IR_REG_4__SCAN_IN,
IR_REG_5__SCAN_IN,
IR_REG_6__SCAN_IN,
IR_REG_7__SCAN_IN,
IR_REG_8__SCAN_IN,
IR_REG_9__SCAN_IN,
IR_REG_10__SCAN_IN,
IR_REG_11__SCAN_IN,
IR_REG_12__SCAN_IN,
IR_REG_13__SCAN_IN,
IR_REG_14__SCAN_IN,
IR_REG_15__SCAN_IN,
IR_REG_16__SCAN_IN,
IR_REG_17__SCAN_IN,
IR_REG_18__SCAN_IN,
IR_REG_19__SCAN_IN,
IR_REG_20__SCAN_IN,
IR_REG_21__SCAN_IN,
IR_REG_22__SCAN_IN,
IR_REG_23__SCAN_IN,
IR_REG_24__SCAN_IN,
IR_REG_25__SCAN_IN,
IR_REG_26__SCAN_IN,
IR_REG_27__SCAN_IN,
IR_REG_28__SCAN_IN,
IR_REG_29__SCAN_IN,
IR_REG_30__SCAN_IN,
IR_REG_31__SCAN_IN,
D_REG_0__SCAN_IN,
D_REG_1__SCAN_IN,
D_REG_2__SCAN_IN,
D_REG_3__SCAN_IN,
D_REG_4__SCAN_IN,
D_REG_5__SCAN_IN,
D_REG_6__SCAN_IN,
D_REG_7__SCAN_IN,
D_REG_8__SCAN_IN,
D_REG_9__SCAN_IN,
D_REG_10__SCAN_IN,
D_REG_11__SCAN_IN,
D_REG_12__SCAN_IN,
D_REG_13__SCAN_IN,
D_REG_14__SCAN_IN,
D_REG_15__SCAN_IN,
D_REG_16__SCAN_IN,
D_REG_17__SCAN_IN,
D_REG_18__SCAN_IN,
D_REG_19__SCAN_IN,
D_REG_20__SCAN_IN,
D_REG_21__SCAN_IN,
D_REG_22__SCAN_IN,
D_REG_23__SCAN_IN,
D_REG_24__SCAN_IN,
D_REG_25__SCAN_IN,
D_REG_26__SCAN_IN,
D_REG_27__SCAN_IN,
D_REG_28__SCAN_IN,
D_REG_29__SCAN_IN,
D_REG_30__SCAN_IN,
D_REG_31__SCAN_IN,
REG0_REG_0__SCAN_IN,
REG0_REG_1__SCAN_IN,
REG0_REG_2__SCAN_IN,
REG0_REG_3__SCAN_IN,
REG0_REG_4__SCAN_IN,
REG0_REG_5__SCAN_IN,
REG0_REG_6__SCAN_IN,
REG0_REG_7__SCAN_IN,
REG0_REG_8__SCAN_IN,
REG0_REG_9__SCAN_IN,
REG0_REG_10__SCAN_IN,
REG0_REG_11__SCAN_IN,
REG0_REG_12__SCAN_IN,
REG0_REG_13__SCAN_IN,
REG0_REG_14__SCAN_IN,
REG0_REG_15__SCAN_IN,
REG0_REG_16__SCAN_IN,
REG0_REG_17__SCAN_IN,
REG0_REG_18__SCAN_IN,
REG0_REG_19__SCAN_IN,
REG0_REG_20__SCAN_IN,
REG0_REG_21__SCAN_IN,
REG0_REG_22__SCAN_IN,
REG0_REG_23__SCAN_IN,
REG0_REG_24__SCAN_IN,
REG0_REG_25__SCAN_IN,
REG0_REG_26__SCAN_IN,
REG0_REG_27__SCAN_IN,
REG0_REG_28__SCAN_IN,
REG0_REG_29__SCAN_IN,
REG0_REG_30__SCAN_IN,
REG0_REG_31__SCAN_IN,
REG1_REG_0__SCAN_IN,
REG1_REG_1__SCAN_IN,
REG1_REG_2__SCAN_IN,
REG1_REG_3__SCAN_IN,
REG1_REG_4__SCAN_IN,
REG1_REG_5__SCAN_IN,
REG1_REG_6__SCAN_IN,
REG1_REG_7__SCAN_IN,
REG1_REG_8__SCAN_IN,
REG1_REG_9__SCAN_IN,
REG1_REG_10__SCAN_IN,
REG1_REG_11__SCAN_IN,
REG1_REG_12__SCAN_IN,
REG1_REG_13__SCAN_IN,
REG1_REG_14__SCAN_IN,
REG1_REG_15__SCAN_IN,
REG1_REG_16__SCAN_IN,
REG1_REG_17__SCAN_IN,
REG1_REG_18__SCAN_IN,
REG1_REG_19__SCAN_IN,
REG1_REG_20__SCAN_IN,
REG1_REG_21__SCAN_IN,
REG1_REG_22__SCAN_IN,
REG1_REG_23__SCAN_IN,
REG1_REG_24__SCAN_IN,
REG1_REG_25__SCAN_IN,
REG1_REG_26__SCAN_IN,
REG1_REG_27__SCAN_IN,
REG1_REG_28__SCAN_IN,
REG1_REG_29__SCAN_IN,
REG1_REG_30__SCAN_IN,
REG1_REG_31__SCAN_IN,
REG2_REG_0__SCAN_IN,
REG2_REG_1__SCAN_IN,
REG2_REG_2__SCAN_IN,
REG2_REG_3__SCAN_IN,
REG2_REG_4__SCAN_IN,
REG2_REG_5__SCAN_IN,
REG2_REG_6__SCAN_IN,
REG2_REG_7__SCAN_IN,
REG2_REG_8__SCAN_IN,
REG2_REG_9__SCAN_IN,
REG2_REG_10__SCAN_IN,
REG2_REG_11__SCAN_IN,
REG2_REG_12__SCAN_IN,
REG2_REG_13__SCAN_IN,
REG2_REG_14__SCAN_IN,
REG2_REG_15__SCAN_IN,
REG2_REG_16__SCAN_IN,
REG2_REG_17__SCAN_IN,
REG2_REG_18__SCAN_IN,
REG2_REG_19__SCAN_IN,
REG2_REG_20__SCAN_IN,
REG2_REG_21__SCAN_IN,
REG2_REG_22__SCAN_IN,
REG2_REG_23__SCAN_IN,
REG2_REG_24__SCAN_IN,
REG2_REG_25__SCAN_IN,
REG2_REG_26__SCAN_IN,
REG2_REG_27__SCAN_IN,
REG2_REG_28__SCAN_IN,
REG2_REG_29__SCAN_IN,
REG2_REG_30__SCAN_IN,
REG2_REG_31__SCAN_IN,
ADDR_REG_19__SCAN_IN,
ADDR_REG_18__SCAN_IN,
ADDR_REG_17__SCAN_IN,
ADDR_REG_16__SCAN_IN,
ADDR_REG_15__SCAN_IN,
ADDR_REG_14__SCAN_IN,
ADDR_REG_13__SCAN_IN,
ADDR_REG_12__SCAN_IN,
ADDR_REG_11__SCAN_IN,
ADDR_REG_10__SCAN_IN,
ADDR_REG_9__SCAN_IN,
ADDR_REG_8__SCAN_IN,
ADDR_REG_7__SCAN_IN,
ADDR_REG_6__SCAN_IN,
ADDR_REG_5__SCAN_IN,
ADDR_REG_4__SCAN_IN,
ADDR_REG_3__SCAN_IN,
ADDR_REG_2__SCAN_IN,
ADDR_REG_1__SCAN_IN,
ADDR_REG_0__SCAN_IN,
DATAO_REG_0__SCAN_IN,
DATAO_REG_1__SCAN_IN,
DATAO_REG_2__SCAN_IN,
DATAO_REG_3__SCAN_IN,
DATAO_REG_4__SCAN_IN,
DATAO_REG_5__SCAN_IN,
DATAO_REG_6__SCAN_IN,
DATAO_REG_7__SCAN_IN,
DATAO_REG_8__SCAN_IN,
DATAO_REG_9__SCAN_IN,
DATAO_REG_10__SCAN_IN,
DATAO_REG_11__SCAN_IN,
DATAO_REG_12__SCAN_IN,
DATAO_REG_13__SCAN_IN,
DATAO_REG_14__SCAN_IN,
DATAO_REG_15__SCAN_IN,
DATAO_REG_16__SCAN_IN,
DATAO_REG_17__SCAN_IN,
DATAO_REG_18__SCAN_IN,
DATAO_REG_19__SCAN_IN,
DATAO_REG_20__SCAN_IN,
DATAO_REG_21__SCAN_IN,
DATAO_REG_22__SCAN_IN,
DATAO_REG_23__SCAN_IN,
DATAO_REG_24__SCAN_IN,
DATAO_REG_25__SCAN_IN,
DATAO_REG_26__SCAN_IN,
DATAO_REG_27__SCAN_IN,
DATAO_REG_28__SCAN_IN,
DATAO_REG_29__SCAN_IN,
DATAO_REG_30__SCAN_IN,
DATAO_REG_31__SCAN_IN,
B_REG_SCAN_IN,
REG3_REG_15__SCAN_IN,
REG3_REG_26__SCAN_IN,
REG3_REG_6__SCAN_IN,
REG3_REG_18__SCAN_IN,
REG3_REG_2__SCAN_IN,
REG3_REG_11__SCAN_IN,
REG3_REG_22__SCAN_IN,
U3352,
U3351,
U3350,
U3349,
U3348,
U3347,
U3346,
U3345,
U3344,
U3343,
U3342,
U3341,
U3340,
U3339,
U3338,
U3337,
U3336,
U3335,
U3334,
U3333,
U3332,
U3331,
U3330,
U3329,
U3328,
U3327,
U3326,
U3325,
U3324,
U3323,
U3322,
U3321,
U3458,
U3459,
U3320,
U3319,
U3318,
U3317,
U3316,
U3315,
U3314,
U3313,
U3312,
U3311,
U3310,
U3309,
U3308,
U3307,
U3306,
U3305,
U3304,
U3303,
U3302,
U3301,
U3300,
U3299,
U3298,
U3297,
U3296,
U3295,
U3294,
U3293,
U3292,
U3291,
U3467,
U3469,
U3471,
U3473,
U3475,
U3477,
U3479,
U3481,
U3483,
U3485,
U3487,
U3489,
U3491,
U3493,
U3495,
U3497,
U3499,
U3501,
U3503,
U3505,
U3506,
U3507,
U3508,
U3509,
U3510,
U3511,
U3512,
U3513,
U3514,
U3515,
U3516,
U3517,
U3518,
U3519,
U3520,
U3521,
U3522,
U3523,
U3524,
U3525,
U3526,
U3527,
U3528,
U3529,
U3530,
U3531,
U3532,
U3533,
U3534,
U3535,
U3536,
U3537,
U3538,
U3539,
U3540,
U3541,
U3542,
U3543,
U3544,
U3545,
U3546,
U3547,
U3548,
U3549,
U3290,
U3289,
U3288,
U3287,
U3286,
U3285,
U3284,
U3283,
U3282,
U3281,
U3280,
U3279,
U3278,
U3277,
U3276,
U3275,
U3274,
U3273,
U3272,
U3271,
U3270,
U3269,
U3268,
U3267,
U3266,
U3265,
U3264,
U3263,
U3262,
U3354,
U3261,
U3260,
U3259,
U3258,
U3257,
U3256,
U3255,
U3254,
U3253,
U3252,
U3251,
U3250,
U3249,
U3248,
U3247,
U3246,
U3245,
U3244,
U3243,
U3242,
U3241,
U3240,
U3550,
U3551,
U3552,
U3553,
U3554,
U3555,
U3556,
U3557,
U3558,
U3559,
U3560,
U3561,
U3562,
U3563,
U3564,
U3565,
U3566,
U3567,
U3568,
U3569,
U3570,
U3571,
U3572,
U3573,
U3574,
U3575,
U3576,
U3577,
U3578,
U3579,
U3580,
U3581,
U3239,
U3238,
U3237,
U3236,
U3235,
U3234,
U3233,
U3232,
U3231,
U3230,
U3229,
U3228,
U3227,
U3226,
U3225,
U3224,
U3223,
U3222,
U3221,
U3220,
U3219,
U3218,
U3217,
U3216,
U3215,
U3214,
U3213,
U3212,
U3211,
U3210,
U3149,
U3148,
U4043);

input DATAI_31_;
input DATAI_30_;
input DATAI_29_;
input DATAI_28_;
input DATAI_27_;
input DATAI_26_;
input DATAI_25_;
input DATAI_24_;
input DATAI_23_;
input DATAI_22_;
input DATAI_21_;
input DATAI_20_;
input DATAI_19_;
input DATAI_18_;
input DATAI_17_;
input DATAI_16_;
input DATAI_15_;
input DATAI_14_;
input DATAI_13_;
input DATAI_12_;
input DATAI_11_;
input DATAI_10_;
input DATAI_9_;
input DATAI_8_;
input DATAI_7_;
input DATAI_6_;
input DATAI_5_;
input DATAI_4_;
input DATAI_3_;
input DATAI_2_;
input DATAI_1_;
input DATAI_0_;
input STATE_REG_SCAN_IN;
input REG3_REG_7__SCAN_IN;
input REG3_REG_27__SCAN_IN;
input REG3_REG_14__SCAN_IN;
input REG3_REG_23__SCAN_IN;
input REG3_REG_10__SCAN_IN;
input REG3_REG_3__SCAN_IN;
input REG3_REG_19__SCAN_IN;
input REG3_REG_28__SCAN_IN;
input REG3_REG_8__SCAN_IN;
input REG3_REG_1__SCAN_IN;
input REG3_REG_21__SCAN_IN;
input REG3_REG_12__SCAN_IN;
input REG3_REG_25__SCAN_IN;
input REG3_REG_16__SCAN_IN;
input REG3_REG_5__SCAN_IN;
input REG3_REG_17__SCAN_IN;
input REG3_REG_24__SCAN_IN;
input REG3_REG_4__SCAN_IN;
input REG3_REG_9__SCAN_IN;
input REG3_REG_0__SCAN_IN;
input REG3_REG_20__SCAN_IN;
input REG3_REG_13__SCAN_IN;
input IR_REG_0__SCAN_IN;
input IR_REG_1__SCAN_IN;
input IR_REG_2__SCAN_IN;
input IR_REG_3__SCAN_IN;
input IR_REG_4__SCAN_IN;
input IR_REG_5__SCAN_IN;
input IR_REG_6__SCAN_IN;
input IR_REG_7__SCAN_IN;
input IR_REG_8__SCAN_IN;
input IR_REG_9__SCAN_IN;
input IR_REG_10__SCAN_IN;
input IR_REG_11__SCAN_IN;
input IR_REG_12__SCAN_IN;
input IR_REG_13__SCAN_IN;
input IR_REG_14__SCAN_IN;
input IR_REG_15__SCAN_IN;
input IR_REG_16__SCAN_IN;
input IR_REG_17__SCAN_IN;
input IR_REG_18__SCAN_IN;
input IR_REG_19__SCAN_IN;
input IR_REG_20__SCAN_IN;
input IR_REG_21__SCAN_IN;
input IR_REG_22__SCAN_IN;
input IR_REG_23__SCAN_IN;
input IR_REG_24__SCAN_IN;
input IR_REG_25__SCAN_IN;
input IR_REG_26__SCAN_IN;
input IR_REG_27__SCAN_IN;
input IR_REG_28__SCAN_IN;
input IR_REG_29__SCAN_IN;
input IR_REG_30__SCAN_IN;
input IR_REG_31__SCAN_IN;
input D_REG_0__SCAN_IN;
input D_REG_1__SCAN_IN;
input D_REG_2__SCAN_IN;
input D_REG_3__SCAN_IN;
input D_REG_4__SCAN_IN;
input D_REG_5__SCAN_IN;
input D_REG_6__SCAN_IN;
input D_REG_7__SCAN_IN;
input D_REG_8__SCAN_IN;
input D_REG_9__SCAN_IN;
input D_REG_10__SCAN_IN;
input D_REG_11__SCAN_IN;
input D_REG_12__SCAN_IN;
input D_REG_13__SCAN_IN;
input D_REG_14__SCAN_IN;
input D_REG_15__SCAN_IN;
input D_REG_16__SCAN_IN;
input D_REG_17__SCAN_IN;
input D_REG_18__SCAN_IN;
input D_REG_19__SCAN_IN;
input D_REG_20__SCAN_IN;
input D_REG_21__SCAN_IN;
input D_REG_22__SCAN_IN;
input D_REG_23__SCAN_IN;
input D_REG_24__SCAN_IN;
input D_REG_25__SCAN_IN;
input D_REG_26__SCAN_IN;
input D_REG_27__SCAN_IN;
input D_REG_28__SCAN_IN;
input D_REG_29__SCAN_IN;
input D_REG_30__SCAN_IN;
input D_REG_31__SCAN_IN;
input REG0_REG_0__SCAN_IN;
input REG0_REG_1__SCAN_IN;
input REG0_REG_2__SCAN_IN;
input REG0_REG_3__SCAN_IN;
input REG0_REG_4__SCAN_IN;
input REG0_REG_5__SCAN_IN;
input REG0_REG_6__SCAN_IN;
input REG0_REG_7__SCAN_IN;
input REG0_REG_8__SCAN_IN;
input REG0_REG_9__SCAN_IN;
input REG0_REG_10__SCAN_IN;
input REG0_REG_11__SCAN_IN;
input REG0_REG_12__SCAN_IN;
input REG0_REG_13__SCAN_IN;
input REG0_REG_14__SCAN_IN;
input REG0_REG_15__SCAN_IN;
input REG0_REG_16__SCAN_IN;
input REG0_REG_17__SCAN_IN;
input REG0_REG_18__SCAN_IN;
input REG0_REG_19__SCAN_IN;
input REG0_REG_20__SCAN_IN;
input REG0_REG_21__SCAN_IN;
input REG0_REG_22__SCAN_IN;
input REG0_REG_23__SCAN_IN;
input REG0_REG_24__SCAN_IN;
input REG0_REG_25__SCAN_IN;
input REG0_REG_26__SCAN_IN;
input REG0_REG_27__SCAN_IN;
input REG0_REG_28__SCAN_IN;
input REG0_REG_29__SCAN_IN;
input REG0_REG_30__SCAN_IN;
input REG0_REG_31__SCAN_IN;
input REG1_REG_0__SCAN_IN;
input REG1_REG_1__SCAN_IN;
input REG1_REG_2__SCAN_IN;
input REG1_REG_3__SCAN_IN;
input REG1_REG_4__SCAN_IN;
input REG1_REG_5__SCAN_IN;
input REG1_REG_6__SCAN_IN;
input REG1_REG_7__SCAN_IN;
input REG1_REG_8__SCAN_IN;
input REG1_REG_9__SCAN_IN;
input REG1_REG_10__SCAN_IN;
input REG1_REG_11__SCAN_IN;
input REG1_REG_12__SCAN_IN;
input REG1_REG_13__SCAN_IN;
input REG1_REG_14__SCAN_IN;
input REG1_REG_15__SCAN_IN;
input REG1_REG_16__SCAN_IN;
input REG1_REG_17__SCAN_IN;
input REG1_REG_18__SCAN_IN;
input REG1_REG_19__SCAN_IN;
input REG1_REG_20__SCAN_IN;
input REG1_REG_21__SCAN_IN;
input REG1_REG_22__SCAN_IN;
input REG1_REG_23__SCAN_IN;
input REG1_REG_24__SCAN_IN;
input REG1_REG_25__SCAN_IN;
input REG1_REG_26__SCAN_IN;
input REG1_REG_27__SCAN_IN;
input REG1_REG_28__SCAN_IN;
input REG1_REG_29__SCAN_IN;
input REG1_REG_30__SCAN_IN;
input REG1_REG_31__SCAN_IN;
input REG2_REG_0__SCAN_IN;
input REG2_REG_1__SCAN_IN;
input REG2_REG_2__SCAN_IN;
input REG2_REG_3__SCAN_IN;
input REG2_REG_4__SCAN_IN;
input REG2_REG_5__SCAN_IN;
input REG2_REG_6__SCAN_IN;
input REG2_REG_7__SCAN_IN;
input REG2_REG_8__SCAN_IN;
input REG2_REG_9__SCAN_IN;
input REG2_REG_10__SCAN_IN;
input REG2_REG_11__SCAN_IN;
input REG2_REG_12__SCAN_IN;
input REG2_REG_13__SCAN_IN;
input REG2_REG_14__SCAN_IN;
input REG2_REG_15__SCAN_IN;
input REG2_REG_16__SCAN_IN;
input REG2_REG_17__SCAN_IN;
input REG2_REG_18__SCAN_IN;
input REG2_REG_19__SCAN_IN;
input REG2_REG_20__SCAN_IN;
input REG2_REG_21__SCAN_IN;
input REG2_REG_22__SCAN_IN;
input REG2_REG_23__SCAN_IN;
input REG2_REG_24__SCAN_IN;
input REG2_REG_25__SCAN_IN;
input REG2_REG_26__SCAN_IN;
input REG2_REG_27__SCAN_IN;
input REG2_REG_28__SCAN_IN;
input REG2_REG_29__SCAN_IN;
input REG2_REG_30__SCAN_IN;
input REG2_REG_31__SCAN_IN;
input ADDR_REG_19__SCAN_IN;
input ADDR_REG_18__SCAN_IN;
input ADDR_REG_17__SCAN_IN;
input ADDR_REG_16__SCAN_IN;
input ADDR_REG_15__SCAN_IN;
input ADDR_REG_14__SCAN_IN;
input ADDR_REG_13__SCAN_IN;
input ADDR_REG_12__SCAN_IN;
input ADDR_REG_11__SCAN_IN;
input ADDR_REG_10__SCAN_IN;
input ADDR_REG_9__SCAN_IN;
input ADDR_REG_8__SCAN_IN;
input ADDR_REG_7__SCAN_IN;
input ADDR_REG_6__SCAN_IN;
input ADDR_REG_5__SCAN_IN;
input ADDR_REG_4__SCAN_IN;
input ADDR_REG_3__SCAN_IN;
input ADDR_REG_2__SCAN_IN;
input ADDR_REG_1__SCAN_IN;
input ADDR_REG_0__SCAN_IN;
input DATAO_REG_0__SCAN_IN;
input DATAO_REG_1__SCAN_IN;
input DATAO_REG_2__SCAN_IN;
input DATAO_REG_3__SCAN_IN;
input DATAO_REG_4__SCAN_IN;
input DATAO_REG_5__SCAN_IN;
input DATAO_REG_6__SCAN_IN;
input DATAO_REG_7__SCAN_IN;
input DATAO_REG_8__SCAN_IN;
input DATAO_REG_9__SCAN_IN;
input DATAO_REG_10__SCAN_IN;
input DATAO_REG_11__SCAN_IN;
input DATAO_REG_12__SCAN_IN;
input DATAO_REG_13__SCAN_IN;
input DATAO_REG_14__SCAN_IN;
input DATAO_REG_15__SCAN_IN;
input DATAO_REG_16__SCAN_IN;
input DATAO_REG_17__SCAN_IN;
input DATAO_REG_18__SCAN_IN;
input DATAO_REG_19__SCAN_IN;
input DATAO_REG_20__SCAN_IN;
input DATAO_REG_21__SCAN_IN;
input DATAO_REG_22__SCAN_IN;
input DATAO_REG_23__SCAN_IN;
input DATAO_REG_24__SCAN_IN;
input DATAO_REG_25__SCAN_IN;
input DATAO_REG_26__SCAN_IN;
input DATAO_REG_27__SCAN_IN;
input DATAO_REG_28__SCAN_IN;
input DATAO_REG_29__SCAN_IN;
input DATAO_REG_30__SCAN_IN;
input DATAO_REG_31__SCAN_IN;
input B_REG_SCAN_IN;
input REG3_REG_15__SCAN_IN;
input REG3_REG_26__SCAN_IN;
input REG3_REG_6__SCAN_IN;
input REG3_REG_18__SCAN_IN;
input REG3_REG_2__SCAN_IN;
input REG3_REG_11__SCAN_IN;
input REG3_REG_22__SCAN_IN;

output U3352;
output U3351;
output U3350;
output U3349;
output U3348;
output U3347;
output U3346;
output U3345;
output U3344;
output U3343;
output U3342;
output U3341;
output U3340;
output U3339;
output U3338;
output U3337;
output U3336;
output U3335;
output U3334;
output U3333;
output U3332;
output U3331;
output U3330;
output U3329;
output U3328;
output U3327;
output U3326;
output U3325;
output U3324;
output U3323;
output U3322;
output U3321;
output U3458;
output U3459;
output U3320;
output U3319;
output U3318;
output U3317;
output U3316;
output U3315;
output U3314;
output U3313;
output U3312;
output U3311;
output U3310;
output U3309;
output U3308;
output U3307;
output U3306;
output U3305;
output U3304;
output U3303;
output U3302;
output U3301;
output U3300;
output U3299;
output U3298;
output U3297;
output U3296;
output U3295;
output U3294;
output U3293;
output U3292;
output U3291;
output U3467;
output U3469;
output U3471;
output U3473;
output U3475;
output U3477;
output U3479;
output U3481;
output U3483;
output U3485;
output U3487;
output U3489;
output U3491;
output U3493;
output U3495;
output U3497;
output U3499;
output U3501;
output U3503;
output U3505;
output U3506;
output U3507;
output U3508;
output U3509;
output U3510;
output U3511;
output U3512;
output U3513;
output U3514;
output U3515;
output U3516;
output U3517;
output U3518;
output U3519;
output U3520;
output U3521;
output U3522;
output U3523;
output U3524;
output U3525;
output U3526;
output U3527;
output U3528;
output U3529;
output U3530;
output U3531;
output U3532;
output U3533;
output U3534;
output U3535;
output U3536;
output U3537;
output U3538;
output U3539;
output U3540;
output U3541;
output U3542;
output U3543;
output U3544;
output U3545;
output U3546;
output U3547;
output U3548;
output U3549;
output U3290;
output U3289;
output U3288;
output U3287;
output U3286;
output U3285;
output U3284;
output U3283;
output U3282;
output U3281;
output U3280;
output U3279;
output U3278;
output U3277;
output U3276;
output U3275;
output U3274;
output U3273;
output U3272;
output U3271;
output U3270;
output U3269;
output U3268;
output U3267;
output U3266;
output U3265;
output U3264;
output U3263;
output U3262;
output U3354;
output U3261;
output U3260;
output U3259;
output U3258;
output U3257;
output U3256;
output U3255;
output U3254;
output U3253;
output U3252;
output U3251;
output U3250;
output U3249;
output U3248;
output U3247;
output U3246;
output U3245;
output U3244;
output U3243;
output U3242;
output U3241;
output U3240;
output U3550;
output U3551;
output U3552;
output U3553;
output U3554;
output U3555;
output U3556;
output U3557;
output U3558;
output U3559;
output U3560;
output U3561;
output U3562;
output U3563;
output U3564;
output U3565;
output U3566;
output U3567;
output U3568;
output U3569;
output U3570;
output U3571;
output U3572;
output U3573;
output U3574;
output U3575;
output U3576;
output U3577;
output U3578;
output U3579;
output U3580;
output U3581;
output U3239;
output U3238;
output U3237;
output U3236;
output U3235;
output U3234;
output U3233;
output U3232;
output U3231;
output U3230;
output U3229;
output U3228;
output U3227;
output U3226;
output U3225;
output U3224;
output U3223;
output U3222;
output U3221;
output U3220;
output U3219;
output U3218;
output U3217;
output U3216;
output U3215;
output U3214;
output U3213;
output U3212;
output U3211;
output U3210;
output U3149;
output U3148;
output U4043;

wire FE_RN_3_0;
wire FE_RN_2_0;
wire FE_OFN27_n11469;
wire FE_OFN23_n11469;
wire FE_OFN22_n12925;
wire FE_OFN21_n13759;
wire FE_RN_0_0;
wire FE_OFN20_n11698;
wire FE_OFN16_n11466;
wire FE_OFN14_n11467;
wire FE_OFN13_n11467;
wire FE_OFN12_n11467;
wire FE_OFN11_n11467;
wire FE_OFN10_n13571;
wire FE_OFN9_n13503;
wire FE_OFN8_n11821;
wire FE_OFN7_n13835;
wire FE_OFN6_n13667;
wire FE_OFN5_n12926;
wire FE_OFN3_n13832;
wire FE_OFN2_n13580;
wire FE_OFN1_n13320;
wire FE_OFN0_n11847;
wire FE_DBTN1_n11467;
wire FE_DBTN0_n11469;
wire n11157;
wire n11159;
wire n11160;
wire n11161;
wire n11164;
wire n11165;
wire n11166;
wire n11167;
wire n11169;
wire n11170;
wire n11171;
wire n11172;
wire n11173;
wire n11174;
wire n11175;
wire n11176;
wire n11177;
wire n11178;
wire n11179;
wire n11181;
wire n11182;
wire n11183;
wire n11184;
wire n11186;
wire n11187;
wire n11189;
wire n11190;
wire n11191;
wire n11192;
wire n11193;
wire n11194;
wire n11195;
wire n11196;
wire n11197;
wire n11201;
wire n11202;
wire n11203;
wire n11204;
wire n11205;
wire n11206;
wire n11207;
wire n11208;
wire n11209;
wire n11210;
wire n11211;
wire n11212;
wire n11213;
wire n11214;
wire n11215;
wire n11216;
wire n11217;
wire n11218;
wire n11219;
wire n11220;
wire n11222;
wire n11223;
wire n11224;
wire n11225;
wire n11226;
wire n11227;
wire n11228;
wire n11229;
wire n11230;
wire n11231;
wire n11232;
wire n11233;
wire n11234;
wire n11235;
wire n11236;
wire n11237;
wire n11238;
wire n11239;
wire n11240;
wire n11241;
wire n11242;
wire n11243;
wire n11244;
wire n11245;
wire n11246;
wire n11247;
wire n11248;
wire n11249;
wire n11250;
wire n11251;
wire n11252;
wire n11253;
wire n11254;
wire n11255;
wire n11256;
wire n11257;
wire n11258;
wire n11259;
wire n11260;
wire n11261;
wire n11262;
wire n11263;
wire n11264;
wire n11265;
wire n11266;
wire n11267;
wire n11268;
wire n11269;
wire n11270;
wire n11271;
wire n11272;
wire n11273;
wire n11274;
wire n11275;
wire n11276;
wire n11277;
wire n11279;
wire n11280;
wire n11282;
wire n11283;
wire n11284;
wire n11286;
wire n11287;
wire n11288;
wire n11289;
wire n11291;
wire n11292;
wire n11293;
wire n11294;
wire n11295;
wire n11296;
wire n11297;
wire n11298;
wire n11299;
wire n11300;
wire n11301;
wire n11303;
wire n11304;
wire n11305;
wire n11306;
wire n11308;
wire n11309;
wire n11310;
wire n11311;
wire n11312;
wire n11313;
wire n11314;
wire n11315;
wire n11316;
wire n11317;
wire n11318;
wire n11319;
wire n11320;
wire n11321;
wire n11322;
wire n11323;
wire n11324;
wire n11325;
wire n11326;
wire n11327;
wire n11328;
wire n11329;
wire n11330;
wire n11332;
wire n11333;
wire n11334;
wire n11335;
wire n11336;
wire n11337;
wire n11340;
wire n11341;
wire n11342;
wire n11343;
wire n11344;
wire n11345;
wire n11346;
wire n11347;
wire n11350;
wire n11351;
wire n11352;
wire n11353;
wire n11354;
wire n11355;
wire n11356;
wire n11357;
wire n11358;
wire n11359;
wire n11360;
wire n11361;
wire n11362;
wire n11363;
wire n11364;
wire n11365;
wire n11366;
wire n11367;
wire n11368;
wire n11369;
wire n11370;
wire n11371;
wire n11372;
wire n11373;
wire n11374;
wire n11375;
wire n11376;
wire n11377;
wire n11378;
wire n11379;
wire n11380;
wire n11381;
wire n11382;
wire n11383;
wire n11384;
wire n11385;
wire n11386;
wire n11387;
wire n11388;
wire n11389;
wire n11390;
wire n11391;
wire n11392;
wire n11393;
wire n11394;
wire n11395;
wire n11396;
wire n11397;
wire n11398;
wire n11399;
wire n11400;
wire n11401;
wire n11402;
wire n11403;
wire n11404;
wire n11405;
wire n11406;
wire n11407;
wire n11408;
wire n11409;
wire n11410;
wire n11411;
wire n11412;
wire n11413;
wire n11414;
wire n11415;
wire n11416;
wire n11417;
wire n11418;
wire n11419;
wire n11420;
wire n11421;
wire n11422;
wire n11423;
wire n11424;
wire n11425;
wire n11426;
wire n11427;
wire n11428;
wire n11429;
wire n11430;
wire n11431;
wire n11432;
wire n11436;
wire n11437;
wire n11438;
wire n11439;
wire n11440;
wire n11441;
wire n11442;
wire n11443;
wire n11444;
wire n11445;
wire n11446;
wire n11447;
wire n11448;
wire n11449;
wire n11450;
wire n11451;
wire n11452;
wire n11454;
wire n11458;
wire n11459;
wire n11460;
wire n11461;
wire n11462;
wire n11463;
wire n11464;
wire n11465;
wire n11466;
wire n11467;
wire n11469;
wire n11470;
wire n11471;
wire n11472;
wire n11473;
wire n11474;
wire n11475;
wire n11476;
wire n11477;
wire n11478;
wire n11479;
wire n11480;
wire n11481;
wire n11482;
wire n11484;
wire n11485;
wire n11486;
wire n11487;
wire n11488;
wire n11489;
wire n11490;
wire n11491;
wire n11492;
wire n11493;
wire n11494;
wire n11495;
wire n11496;
wire n11497;
wire n11498;
wire n11499;
wire n11501;
wire n11502;
wire n11503;
wire n11504;
wire n11505;
wire n11506;
wire n11507;
wire n11508;
wire n11509;
wire n11510;
wire n11511;
wire n11512;
wire n11513;
wire n11514;
wire n11515;
wire n11516;
wire n11517;
wire n11518;
wire n11519;
wire n11520;
wire n11521;
wire n11522;
wire n11523;
wire n11524;
wire n11525;
wire n11526;
wire n11528;
wire n11529;
wire n11530;
wire n11531;
wire n11532;
wire n11533;
wire n11536;
wire n11537;
wire n11538;
wire n11539;
wire n11540;
wire n11541;
wire n11542;
wire n11543;
wire n11544;
wire n11545;
wire n11546;
wire n11547;
wire n11548;
wire n11549;
wire n11550;
wire n11551;
wire n11552;
wire n11553;
wire n11554;
wire n11555;
wire n11556;
wire n11557;
wire n11558;
wire n11559;
wire n11560;
wire n11561;
wire n11562;
wire n11563;
wire n11564;
wire n11567;
wire n11568;
wire n11569;
wire n11571;
wire n11572;
wire n11573;
wire n11574;
wire n11575;
wire n11576;
wire n11577;
wire n11580;
wire n11581;
wire n11582;
wire n11583;
wire n11584;
wire n11585;
wire n11586;
wire n11587;
wire n11590;
wire n11591;
wire n11592;
wire n11593;
wire n11594;
wire n11595;
wire n11596;
wire n11599;
wire n11600;
wire n11601;
wire n11602;
wire n11603;
wire n11604;
wire n11605;
wire n11608;
wire n11609;
wire n11610;
wire n11611;
wire n11612;
wire n11613;
wire n11614;
wire n11615;
wire n11616;
wire n11617;
wire n11618;
wire n11619;
wire n11620;
wire n11621;
wire n11622;
wire n11623;
wire n11624;
wire n11625;
wire n11626;
wire n11627;
wire n11630;
wire n11631;
wire n11632;
wire n11633;
wire n11634;
wire n11635;
wire n11636;
wire n11640;
wire n11641;
wire n11642;
wire n11644;
wire n11645;
wire n11646;
wire n11647;
wire n11648;
wire n11653;
wire n11654;
wire n11655;
wire n11657;
wire n11658;
wire n11660;
wire n11661;
wire n11662;
wire n11664;
wire n11665;
wire n11666;
wire n11667;
wire n11670;
wire n11671;
wire n11672;
wire n11673;
wire n11674;
wire n11675;
wire n11676;
wire n11678;
wire n11679;
wire n11680;
wire n11681;
wire n11682;
wire n11683;
wire n11684;
wire n11685;
wire n11686;
wire n11687;
wire n11689;
wire n11690;
wire n11691;
wire n11692;
wire n11693;
wire n11694;
wire n11695;
wire n11696;
wire n11697;
wire n11698;
wire n11699;
wire n11700;
wire n11701;
wire n11702;
wire n11703;
wire n11704;
wire n11705;
wire n11706;
wire n11707;
wire n11708;
wire n11709;
wire n11710;
wire n11711;
wire n11712;
wire n11713;
wire n11714;
wire n11715;
wire n11716;
wire n11718;
wire n11719;
wire n11720;
wire n11721;
wire n11722;
wire n11723;
wire n11724;
wire n11725;
wire n11726;
wire n11727;
wire n11728;
wire n11729;
wire n11730;
wire n11731;
wire n11732;
wire n11733;
wire n11734;
wire n11735;
wire n11736;
wire n11737;
wire n11738;
wire n11739;
wire n11740;
wire n11741;
wire n11742;
wire n11743;
wire n11744;
wire n11745;
wire n11746;
wire n11747;
wire n11748;
wire n11749;
wire n11750;
wire n11751;
wire n11752;
wire n11753;
wire n11754;
wire n11755;
wire n11756;
wire n11757;
wire n11758;
wire n11759;
wire n11760;
wire n11761;
wire n11764;
wire n11765;
wire n11767;
wire n11768;
wire n11769;
wire n11770;
wire n11772;
wire n11773;
wire n11774;
wire n11775;
wire n11776;
wire n11778;
wire n11779;
wire n11780;
wire n11781;
wire n11782;
wire n11783;
wire n11784;
wire n11785;
wire n11786;
wire n11787;
wire n11789;
wire n11791;
wire n11792;
wire n11794;
wire n11795;
wire n11796;
wire n11797;
wire n11798;
wire n11799;
wire n11800;
wire n11801;
wire n11802;
wire n11803;
wire n11804;
wire n11806;
wire n11807;
wire n11808;
wire n11809;
wire n11810;
wire n11811;
wire n11812;
wire n11815;
wire n11816;
wire n11817;
wire n11818;
wire n11819;
wire n11821;
wire n11822;
wire n11823;
wire n11824;
wire n11825;
wire n11826;
wire n11827;
wire n11828;
wire n11829;
wire n11830;
wire n11831;
wire n11832;
wire n11833;
wire n11834;
wire n11835;
wire n11836;
wire n11837;
wire n11838;
wire n11839;
wire n11840;
wire n11841;
wire n11842;
wire n11843;
wire n11844;
wire n11845;
wire n11846;
wire n11847;
wire n11848;
wire n11849;
wire n11850;
wire n11851;
wire n11852;
wire n11853;
wire n11854;
wire n11855;
wire n11856;
wire n11857;
wire n11858;
wire n11859;
wire n11860;
wire n11861;
wire n11862;
wire n11863;
wire n11864;
wire n11865;
wire n11866;
wire n11867;
wire n11868;
wire n11869;
wire n11870;
wire n11871;
wire n11872;
wire n11873;
wire n11874;
wire n11875;
wire n11876;
wire n11877;
wire n11878;
wire n11879;
wire n11880;
wire n11881;
wire n11882;
wire n11883;
wire n11884;
wire n11885;
wire n11886;
wire n11887;
wire n11888;
wire n11889;
wire n11890;
wire n11891;
wire n11892;
wire n11893;
wire n11894;
wire n11895;
wire n11896;
wire n11900;
wire n11901;
wire n11902;
wire n11903;
wire n11904;
wire n11905;
wire n11906;
wire n11907;
wire n11908;
wire n11909;
wire n11910;
wire n11911;
wire n11912;
wire n11913;
wire n11914;
wire n11915;
wire n11916;
wire n11917;
wire n11918;
wire n11919;
wire n11920;
wire n11921;
wire n11922;
wire n11923;
wire n11924;
wire n11925;
wire n11926;
wire n11927;
wire n11928;
wire n11929;
wire n11930;
wire n11931;
wire n11932;
wire n11933;
wire n11934;
wire n11935;
wire n11938;
wire n11939;
wire n11940;
wire n11941;
wire n11942;
wire n11944;
wire n11945;
wire n11946;
wire n11947;
wire n11948;
wire n11950;
wire n11953;
wire n11954;
wire n11955;
wire n11956;
wire n11957;
wire n11958;
wire n11960;
wire n11961;
wire n11962;
wire n11963;
wire n11964;
wire n11965;
wire n11966;
wire n11967;
wire n11968;
wire n11969;
wire n11970;
wire n11971;
wire n11972;
wire n11973;
wire n11974;
wire n11975;
wire n11976;
wire n11977;
wire n11978;
wire n11979;
wire n11980;
wire n11981;
wire n11982;
wire n11983;
wire n11984;
wire n11985;
wire n11986;
wire n11987;
wire n11988;
wire n11989;
wire n11990;
wire n11991;
wire n11992;
wire n11993;
wire n11994;
wire n11995;
wire n11996;
wire n11997;
wire n11998;
wire n11999;
wire n12000;
wire n12001;
wire n12002;
wire n12003;
wire n12004;
wire n12005;
wire n12006;
wire n12007;
wire n12008;
wire n12009;
wire n12010;
wire n12011;
wire n12012;
wire n12015;
wire n12016;
wire n12019;
wire n12020;
wire n12021;
wire n12022;
wire n12023;
wire n12024;
wire n12025;
wire n12026;
wire n12027;
wire n12028;
wire n12029;
wire n12030;
wire n12031;
wire n12032;
wire n12033;
wire n12034;
wire n12035;
wire n12036;
wire n12037;
wire n12038;
wire n12039;
wire n12040;
wire n12041;
wire n12042;
wire n12045;
wire n12046;
wire n12047;
wire n12048;
wire n12049;
wire n12050;
wire n12051;
wire n12052;
wire n12053;
wire n12054;
wire n12055;
wire n12056;
wire n12057;
wire n12058;
wire n12059;
wire n12060;
wire n12062;
wire n12063;
wire n12064;
wire n12065;
wire n12066;
wire n12067;
wire n12070;
wire n12071;
wire n12072;
wire n12073;
wire n12074;
wire n12075;
wire n12077;
wire n12078;
wire n12079;
wire n12080;
wire n12081;
wire n12084;
wire n12085;
wire n12086;
wire n12087;
wire n12088;
wire n12089;
wire n12090;
wire n12091;
wire n12093;
wire n12094;
wire n12095;
wire n12096;
wire n12097;
wire n12098;
wire n12099;
wire n12100;
wire n12101;
wire n12102;
wire n12103;
wire n12104;
wire n12106;
wire n12107;
wire n12108;
wire n12109;
wire n12110;
wire n12111;
wire n12112;
wire n12113;
wire n12114;
wire n12115;
wire n12116;
wire n12117;
wire n12118;
wire n12119;
wire n12120;
wire n12121;
wire n12124;
wire n12125;
wire n12126;
wire n12127;
wire n12128;
wire n12129;
wire n12130;
wire n12131;
wire n12132;
wire n12133;
wire n12134;
wire n12135;
wire n12136;
wire n12137;
wire n12138;
wire n12139;
wire n12140;
wire n12141;
wire n12142;
wire n12143;
wire n12144;
wire n12145;
wire n12148;
wire n12149;
wire n12150;
wire n12151;
wire n12152;
wire n12155;
wire n12156;
wire n12157;
wire n12158;
wire n12159;
wire n12160;
wire n12161;
wire n12162;
wire n12163;
wire n12164;
wire n12165;
wire n12166;
wire n12167;
wire n12168;
wire n12169;
wire n12170;
wire n12171;
wire n12172;
wire n12174;
wire n12175;
wire n12178;
wire n12179;
wire n12181;
wire n12182;
wire n12183;
wire n12184;
wire n12185;
wire n12186;
wire n12187;
wire n12188;
wire n12189;
wire n12190;
wire n12191;
wire n12192;
wire n12193;
wire n12194;
wire n12195;
wire n12196;
wire n12197;
wire n12198;
wire n12199;
wire n12200;
wire n12201;
wire n12202;
wire n12203;
wire n12204;
wire n12205;
wire n12206;
wire n12207;
wire n12208;
wire n12209;
wire n12210;
wire n12211;
wire n12212;
wire n12213;
wire n12214;
wire n12215;
wire n12216;
wire n12217;
wire n12218;
wire n12219;
wire n12220;
wire n12221;
wire n12222;
wire n12223;
wire n12224;
wire n12225;
wire n12226;
wire n12227;
wire n12228;
wire n12229;
wire n12230;
wire n12231;
wire n12232;
wire n12233;
wire n12234;
wire n12235;
wire n12236;
wire n12237;
wire n12238;
wire n12239;
wire n12240;
wire n12241;
wire n12242;
wire n12243;
wire n12246;
wire n12247;
wire n12248;
wire n12249;
wire n12250;
wire n12251;
wire n12252;
wire n12253;
wire n12254;
wire n12255;
wire n12256;
wire n12257;
wire n12258;
wire n12259;
wire n12260;
wire n12261;
wire n12262;
wire n12263;
wire n12264;
wire n12265;
wire n12266;
wire n12267;
wire n12268;
wire n12269;
wire n12270;
wire n12271;
wire n12272;
wire n12273;
wire n12274;
wire n12275;
wire n12276;
wire n12277;
wire n12278;
wire n12279;
wire n12280;
wire n12281;
wire n12282;
wire n12283;
wire n12284;
wire n12285;
wire n12286;
wire n12287;
wire n12288;
wire n12289;
wire n12290;
wire n12291;
wire n12292;
wire n12293;
wire n12294;
wire n12295;
wire n12296;
wire n12297;
wire n12298;
wire n12299;
wire n12300;
wire n12301;
wire n12302;
wire n12303;
wire n12304;
wire n12305;
wire n12306;
wire n12307;
wire n12308;
wire n12309;
wire n12310;
wire n12311;
wire n12312;
wire n12313;
wire n12314;
wire n12315;
wire n12316;
wire n12317;
wire n12318;
wire n12319;
wire n12320;
wire n12323;
wire n12324;
wire n12325;
wire n12328;
wire n12329;
wire n12330;
wire n12333;
wire n12334;
wire n12337;
wire n12338;
wire n12339;
wire n12340;
wire n12341;
wire n12342;
wire n12343;
wire n12344;
wire n12345;
wire n12346;
wire n12347;
wire n12348;
wire n12349;
wire n12350;
wire n12351;
wire n12352;
wire n12353;
wire n12354;
wire n12355;
wire n12356;
wire n12357;
wire n12358;
wire n12359;
wire n12360;
wire n12361;
wire n12362;
wire n12363;
wire n12364;
wire n12365;
wire n12366;
wire n12367;
wire n12368;
wire n12369;
wire n12370;
wire n12371;
wire n12372;
wire n12373;
wire n12374;
wire n12375;
wire n12376;
wire n12377;
wire n12378;
wire n12379;
wire n12380;
wire n12381;
wire n12382;
wire n12383;
wire n12384;
wire n12385;
wire n12386;
wire n12387;
wire n12388;
wire n12389;
wire n12390;
wire n12391;
wire n12392;
wire n12393;
wire n12394;
wire n12395;
wire n12396;
wire n12397;
wire n12398;
wire n12399;
wire n12400;
wire n12403;
wire n12404;
wire n12405;
wire n12406;
wire n12407;
wire n12408;
wire n12409;
wire n12410;
wire n12411;
wire n12412;
wire n12413;
wire n12414;
wire n12415;
wire n12416;
wire n12417;
wire n12418;
wire n12419;
wire n12420;
wire n12421;
wire n12422;
wire n12423;
wire n12424;
wire n12425;
wire n12426;
wire n12427;
wire n12428;
wire n12429;
wire n12430;
wire n12431;
wire n12432;
wire n12433;
wire n12434;
wire n12435;
wire n12436;
wire n12437;
wire n12438;
wire n12439;
wire n12441;
wire n12442;
wire n12443;
wire n12444;
wire n12446;
wire n12447;
wire n12448;
wire n12449;
wire n12450;
wire n12451;
wire n12452;
wire n12453;
wire n12454;
wire n12455;
wire n12456;
wire n12457;
wire n12458;
wire n12459;
wire n12460;
wire n12461;
wire n12462;
wire n12463;
wire n12464;
wire n12465;
wire n12466;
wire n12467;
wire n12468;
wire n12469;
wire n12470;
wire n12471;
wire n12472;
wire n12473;
wire n12474;
wire n12475;
wire n12476;
wire n12477;
wire n12478;
wire n12479;
wire n12480;
wire n12481;
wire n12482;
wire n12483;
wire n12484;
wire n12485;
wire n12486;
wire n12487;
wire n12488;
wire n12489;
wire n12490;
wire n12491;
wire n12492;
wire n12493;
wire n12494;
wire n12495;
wire n12496;
wire n12497;
wire n12498;
wire n12499;
wire n12500;
wire n12501;
wire n12502;
wire n12503;
wire n12504;
wire n12505;
wire n12506;
wire n12507;
wire n12508;
wire n12509;
wire n12510;
wire n12511;
wire n12512;
wire n12513;
wire n12514;
wire n12515;
wire n12516;
wire n12517;
wire n12518;
wire n12520;
wire n12521;
wire n12522;
wire n12523;
wire n12524;
wire n12525;
wire n12526;
wire n12528;
wire n12529;
wire n12530;
wire n12531;
wire n12532;
wire n12533;
wire n12534;
wire n12535;
wire n12536;
wire n12537;
wire n12538;
wire n12539;
wire n12540;
wire n12541;
wire n12542;
wire n12543;
wire n12544;
wire n12545;
wire n12546;
wire n12547;
wire n12548;
wire n12549;
wire n12550;
wire n12551;
wire n12552;
wire n12553;
wire n12554;
wire n12555;
wire n12556;
wire n12561;
wire n12563;
wire n12564;
wire n12565;
wire n12566;
wire n12567;
wire n12568;
wire n12569;
wire n12570;
wire n12571;
wire n12572;
wire n12573;
wire n12574;
wire n12575;
wire n12576;
wire n12577;
wire n12578;
wire n12579;
wire n12580;
wire n12581;
wire n12582;
wire n12584;
wire n12585;
wire n12586;
wire n12587;
wire n12588;
wire n12589;
wire n12590;
wire n12592;
wire n12593;
wire n12594;
wire n12595;
wire n12596;
wire n12597;
wire n12598;
wire n12599;
wire n12600;
wire n12601;
wire n12603;
wire n12604;
wire n12605;
wire n12606;
wire n12607;
wire n12608;
wire n12609;
wire n12610;
wire n12611;
wire n12612;
wire n12613;
wire n12614;
wire n12615;
wire n12616;
wire n12617;
wire n12618;
wire n12619;
wire n12620;
wire n12621;
wire n12622;
wire n12623;
wire n12624;
wire n12625;
wire n12626;
wire n12627;
wire n12628;
wire n12629;
wire n12630;
wire n12631;
wire n12632;
wire n12633;
wire n12634;
wire n12635;
wire n12636;
wire n12637;
wire n12638;
wire n12639;
wire n12640;
wire n12641;
wire n12642;
wire n12643;
wire n12644;
wire n12645;
wire n12646;
wire n12647;
wire n12648;
wire n12649;
wire n12650;
wire n12651;
wire n12652;
wire n12653;
wire n12654;
wire n12655;
wire n12656;
wire n12657;
wire n12658;
wire n12659;
wire n12660;
wire n12661;
wire n12662;
wire n12663;
wire n12664;
wire n12665;
wire n12666;
wire n12667;
wire n12668;
wire n12669;
wire n12670;
wire n12671;
wire n12672;
wire n12673;
wire n12674;
wire n12675;
wire n12676;
wire n12677;
wire n12678;
wire n12679;
wire n12680;
wire n12681;
wire n12682;
wire n12683;
wire n12684;
wire n12685;
wire n12686;
wire n12687;
wire n12688;
wire n12689;
wire n12690;
wire n12691;
wire n12692;
wire n12693;
wire n12694;
wire n12695;
wire n12696;
wire n12697;
wire n12698;
wire n12699;
wire n12700;
wire n12701;
wire n12702;
wire n12703;
wire n12704;
wire n12705;
wire n12706;
wire n12707;
wire n12708;
wire n12709;
wire n12710;
wire n12711;
wire n12712;
wire n12713;
wire n12714;
wire n12715;
wire n12716;
wire n12717;
wire n12718;
wire n12719;
wire n12720;
wire n12721;
wire n12722;
wire n12723;
wire n12724;
wire n12725;
wire n12726;
wire n12727;
wire n12728;
wire n12729;
wire n12730;
wire n12731;
wire n12732;
wire n12733;
wire n12734;
wire n12735;
wire n12736;
wire n12737;
wire n12738;
wire n12739;
wire n12740;
wire n12741;
wire n12742;
wire n12743;
wire n12744;
wire n12745;
wire n12746;
wire n12747;
wire n12748;
wire n12749;
wire n12750;
wire n12751;
wire n12752;
wire n12753;
wire n12754;
wire n12755;
wire n12756;
wire n12757;
wire n12758;
wire n12759;
wire n12760;
wire n12761;
wire n12762;
wire n12763;
wire n12764;
wire n12765;
wire n12766;
wire n12767;
wire n12768;
wire n12769;
wire n12770;
wire n12771;
wire n12772;
wire n12773;
wire n12774;
wire n12775;
wire n12776;
wire n12778;
wire n12779;
wire n12780;
wire n12781;
wire n12782;
wire n12783;
wire n12784;
wire n12785;
wire n12786;
wire n12787;
wire n12788;
wire n12789;
wire n12790;
wire n12791;
wire n12792;
wire n12793;
wire n12794;
wire n12795;
wire n12796;
wire n12797;
wire n12798;
wire n12799;
wire n12800;
wire n12801;
wire n12802;
wire n12803;
wire n12804;
wire n12805;
wire n12806;
wire n12807;
wire n12808;
wire n12809;
wire n12810;
wire n12811;
wire n12812;
wire n12813;
wire n12815;
wire n12816;
wire n12817;
wire n12818;
wire n12819;
wire n12820;
wire n12821;
wire n12822;
wire n12823;
wire n12824;
wire n12825;
wire n12826;
wire n12827;
wire n12828;
wire n12829;
wire n12830;
wire n12831;
wire n12832;
wire n12833;
wire n12834;
wire n12835;
wire n12836;
wire n12837;
wire n12838;
wire n12839;
wire n12840;
wire n12841;
wire n12843;
wire n12844;
wire n12845;
wire n12846;
wire n12847;
wire n12848;
wire n12849;
wire n12850;
wire n12851;
wire n12852;
wire n12853;
wire n12854;
wire n12855;
wire n12856;
wire n12857;
wire n12858;
wire n12859;
wire n12860;
wire n12861;
wire n12862;
wire n12863;
wire n12864;
wire n12866;
wire n12867;
wire n12868;
wire n12869;
wire n12870;
wire n12871;
wire n12872;
wire n12873;
wire n12874;
wire n12875;
wire n12876;
wire n12877;
wire n12878;
wire n12879;
wire n12880;
wire n12881;
wire n12882;
wire n12883;
wire n12884;
wire n12885;
wire n12886;
wire n12887;
wire n12888;
wire n12889;
wire n12890;
wire n12891;
wire n12892;
wire n12893;
wire n12894;
wire n12895;
wire n12896;
wire n12897;
wire n12898;
wire n12899;
wire n12900;
wire n12901;
wire n12902;
wire n12903;
wire n12904;
wire n12905;
wire n12906;
wire n12907;
wire n12908;
wire n12909;
wire n12910;
wire n12911;
wire n12912;
wire n12913;
wire n12914;
wire n12915;
wire n12916;
wire n12917;
wire n12918;
wire n12919;
wire n12920;
wire n12921;
wire n12922;
wire n12923;
wire n12924;
wire n12925;
wire n12926;
wire n12927;
wire n12928;
wire n12929;
wire n12930;
wire n12931;
wire n12932;
wire n12933;
wire n12934;
wire n12935;
wire n12936;
wire n12937;
wire n12938;
wire n12939;
wire n12940;
wire n12941;
wire n12942;
wire n12943;
wire n12944;
wire n12945;
wire n12947;
wire n12948;
wire n12949;
wire n12950;
wire n12951;
wire n12952;
wire n12953;
wire n12954;
wire n12955;
wire n12956;
wire n12957;
wire n12958;
wire n12959;
wire n12960;
wire n12961;
wire n12962;
wire n12963;
wire n12964;
wire n12965;
wire n12966;
wire n12967;
wire n12968;
wire n12969;
wire n12970;
wire n12971;
wire n12972;
wire n12973;
wire n12974;
wire n12975;
wire n12976;
wire n12977;
wire n12978;
wire n12979;
wire n12980;
wire n12981;
wire n12982;
wire n12983;
wire n12984;
wire n12985;
wire n12986;
wire n12987;
wire n12988;
wire n12989;
wire n12990;
wire n12991;
wire n12992;
wire n12993;
wire n12994;
wire n12995;
wire n12996;
wire n12997;
wire n12998;
wire n12999;
wire n13000;
wire n13001;
wire n13002;
wire n13003;
wire n13004;
wire n13005;
wire n13006;
wire n13007;
wire n13008;
wire n13009;
wire n13010;
wire n13011;
wire n13012;
wire n13013;
wire n13014;
wire n13015;
wire n13016;
wire n13017;
wire n13018;
wire n13019;
wire n13020;
wire n13021;
wire n13022;
wire n13023;
wire n13024;
wire n13025;
wire n13026;
wire n13027;
wire n13028;
wire n13029;
wire n13030;
wire n13031;
wire n13032;
wire n13033;
wire n13034;
wire n13035;
wire n13036;
wire n13037;
wire n13038;
wire n13039;
wire n13040;
wire n13041;
wire n13042;
wire n13043;
wire n13044;
wire n13045;
wire n13048;
wire n13049;
wire n13050;
wire n13051;
wire n13052;
wire n13053;
wire n13054;
wire n13055;
wire n13056;
wire n13057;
wire n13058;
wire n13059;
wire n13060;
wire n13061;
wire n13062;
wire n13063;
wire n13064;
wire n13065;
wire n13066;
wire n13067;
wire n13068;
wire n13069;
wire n13070;
wire n13071;
wire n13072;
wire n13073;
wire n13074;
wire n13075;
wire n13076;
wire n13077;
wire n13078;
wire n13079;
wire n13080;
wire n13081;
wire n13082;
wire n13083;
wire n13084;
wire n13085;
wire n13086;
wire n13087;
wire n13088;
wire n13089;
wire n13090;
wire n13091;
wire n13092;
wire n13093;
wire n13094;
wire n13095;
wire n13096;
wire n13097;
wire n13098;
wire n13099;
wire n13100;
wire n13101;
wire n13102;
wire n13104;
wire n13105;
wire n13106;
wire n13107;
wire n13108;
wire n13109;
wire n13110;
wire n13111;
wire n13112;
wire n13113;
wire n13114;
wire n13115;
wire n13116;
wire n13117;
wire n13118;
wire n13119;
wire n13120;
wire n13121;
wire n13122;
wire n13123;
wire n13124;
wire n13125;
wire n13126;
wire n13127;
wire n13128;
wire n13129;
wire n13130;
wire n13131;
wire n13132;
wire n13133;
wire n13134;
wire n13135;
wire n13136;
wire n13137;
wire n13138;
wire n13139;
wire n13141;
wire n13142;
wire n13143;
wire n13144;
wire n13145;
wire n13146;
wire n13147;
wire n13148;
wire n13149;
wire n13150;
wire n13151;
wire n13152;
wire n13153;
wire n13154;
wire n13155;
wire n13156;
wire n13157;
wire n13158;
wire n13159;
wire n13160;
wire n13161;
wire n13162;
wire n13163;
wire n13164;
wire n13165;
wire n13166;
wire n13167;
wire n13168;
wire n13169;
wire n13170;
wire n13171;
wire n13172;
wire n13173;
wire n13174;
wire n13175;
wire n13176;
wire n13177;
wire n13178;
wire n13179;
wire n13180;
wire n13181;
wire n13182;
wire n13183;
wire n13184;
wire n13185;
wire n13186;
wire n13187;
wire n13188;
wire n13189;
wire n13190;
wire n13191;
wire n13192;
wire n13193;
wire n13194;
wire n13195;
wire n13196;
wire n13197;
wire n13198;
wire n13199;
wire n13200;
wire n13201;
wire n13202;
wire n13203;
wire n13204;
wire n13205;
wire n13206;
wire n13207;
wire n13208;
wire n13209;
wire n13210;
wire n13211;
wire n13212;
wire n13213;
wire n13214;
wire n13215;
wire n13216;
wire n13217;
wire n13218;
wire n13219;
wire n13220;
wire n13221;
wire n13223;
wire n13225;
wire n13226;
wire n13227;
wire n13228;
wire n13229;
wire n13230;
wire n13231;
wire n13232;
wire n13233;
wire n13234;
wire n13235;
wire n13236;
wire n13237;
wire n13238;
wire n13239;
wire n13240;
wire n13241;
wire n13242;
wire n13243;
wire n13244;
wire n13245;
wire n13246;
wire n13247;
wire n13248;
wire n13249;
wire n13250;
wire n13251;
wire n13252;
wire n13253;
wire n13254;
wire n13255;
wire n13256;
wire n13257;
wire n13258;
wire n13259;
wire n13260;
wire n13261;
wire n13262;
wire n13263;
wire n13264;
wire n13265;
wire n13266;
wire n13267;
wire n13268;
wire n13269;
wire n13270;
wire n13271;
wire n13272;
wire n13273;
wire n13274;
wire n13275;
wire n13278;
wire n13279;
wire n13280;
wire n13283;
wire n13284;
wire n13285;
wire n13286;
wire n13287;
wire n13288;
wire n13289;
wire n13290;
wire n13291;
wire n13292;
wire n13293;
wire n13294;
wire n13295;
wire n13296;
wire n13297;
wire n13298;
wire n13299;
wire n13300;
wire n13301;
wire n13302;
wire n13305;
wire n13306;
wire n13307;
wire n13308;
wire n13309;
wire n13311;
wire n13312;
wire n13313;
wire n13314;
wire n13315;
wire n13316;
wire n13317;
wire n13318;
wire n13319;
wire n13320;
wire n13321;
wire n13322;
wire n13323;
wire n13324;
wire n13325;
wire n13326;
wire n13327;
wire n13328;
wire n13329;
wire n13330;
wire n13331;
wire n13332;
wire n13333;
wire n13334;
wire n13335;
wire n13336;
wire n13337;
wire n13338;
wire n13339;
wire n13340;
wire n13341;
wire n13342;
wire n13343;
wire n13344;
wire n13345;
wire n13346;
wire n13347;
wire n13348;
wire n13349;
wire n13350;
wire n13353;
wire n13354;
wire n13355;
wire n13356;
wire n13357;
wire n13358;
wire n13360;
wire n13361;
wire n13362;
wire n13363;
wire n13364;
wire n13366;
wire n13368;
wire n13369;
wire n13370;
wire n13371;
wire n13372;
wire n13373;
wire n13374;
wire n13375;
wire n13376;
wire n13377;
wire n13378;
wire n13379;
wire n13380;
wire n13381;
wire n13382;
wire n13383;
wire n13384;
wire n13385;
wire n13386;
wire n13387;
wire n13388;
wire n13389;
wire n13390;
wire n13391;
wire n13392;
wire n13393;
wire n13395;
wire n13396;
wire n13397;
wire n13398;
wire n13399;
wire n13400;
wire n13401;
wire n13402;
wire n13403;
wire n13404;
wire n13406;
wire n13407;
wire n13408;
wire n13409;
wire n13410;
wire n13411;
wire n13412;
wire n13413;
wire n13414;
wire n13415;
wire n13416;
wire n13417;
wire n13418;
wire n13419;
wire n13420;
wire n13421;
wire n13422;
wire n13423;
wire n13424;
wire n13426;
wire n13427;
wire n13428;
wire n13430;
wire n13431;
wire n13432;
wire n13433;
wire n13434;
wire n13435;
wire n13436;
wire n13437;
wire n13438;
wire n13439;
wire n13440;
wire n13441;
wire n13442;
wire n13443;
wire n13444;
wire n13445;
wire n13446;
wire n13447;
wire n13448;
wire n13452;
wire n13453;
wire n13454;
wire n13455;
wire n13456;
wire n13457;
wire n13458;
wire n13459;
wire n13460;
wire n13461;
wire n13462;
wire n13463;
wire n13464;
wire n13465;
wire n13466;
wire n13467;
wire n13468;
wire n13469;
wire n13470;
wire n13471;
wire n13472;
wire n13473;
wire n13474;
wire n13475;
wire n13476;
wire n13477;
wire n13478;
wire n13479;
wire n13480;
wire n13481;
wire n13482;
wire n13483;
wire n13484;
wire n13485;
wire n13486;
wire n13487;
wire n13488;
wire n13489;
wire n13490;
wire n13491;
wire n13492;
wire n13493;
wire n13494;
wire n13495;
wire n13496;
wire n13497;
wire n13498;
wire n13499;
wire n13500;
wire n13501;
wire n13502;
wire n13503;
wire n13504;
wire n13505;
wire n13506;
wire n13507;
wire n13508;
wire n13509;
wire n13510;
wire n13511;
wire n13512;
wire n13513;
wire n13514;
wire n13515;
wire n13516;
wire n13517;
wire n13518;
wire n13519;
wire n13520;
wire n13521;
wire n13522;
wire n13523;
wire n13524;
wire n13525;
wire n13526;
wire n13527;
wire n13528;
wire n13529;
wire n13530;
wire n13531;
wire n13533;
wire n13534;
wire n13535;
wire n13536;
wire n13537;
wire n13538;
wire n13539;
wire n13540;
wire n13541;
wire n13542;
wire n13543;
wire n13544;
wire n13545;
wire n13546;
wire n13547;
wire n13548;
wire n13549;
wire n13550;
wire n13551;
wire n13552;
wire n13553;
wire n13554;
wire n13555;
wire n13556;
wire n13557;
wire n13558;
wire n13559;
wire n13561;
wire n13562;
wire n13563;
wire n13564;
wire n13565;
wire n13566;
wire n13567;
wire n13568;
wire n13569;
wire n13570;
wire n13571;
wire n13572;
wire n13573;
wire n13574;
wire n13575;
wire n13576;
wire n13577;
wire n13578;
wire n13579;
wire n13580;
wire n13581;
wire n13582;
wire n13583;
wire n13584;
wire n13585;
wire n13586;
wire n13587;
wire n13588;
wire n13589;
wire n13591;
wire n13592;
wire n13593;
wire n13594;
wire n13595;
wire n13596;
wire n13598;
wire n13600;
wire n13601;
wire n13602;
wire n13603;
wire n13604;
wire n13605;
wire n13606;
wire n13607;
wire n13608;
wire n13609;
wire n13610;
wire n13611;
wire n13612;
wire n13613;
wire n13614;
wire n13615;
wire n13616;
wire n13617;
wire n13618;
wire n13619;
wire n13620;
wire n13621;
wire n13622;
wire n13623;
wire n13624;
wire n13625;
wire n13626;
wire n13627;
wire n13628;
wire n13629;
wire n13630;
wire n13631;
wire n13632;
wire n13633;
wire n13634;
wire n13635;
wire n13636;
wire n13637;
wire n13638;
wire n13639;
wire n13640;
wire n13641;
wire n13642;
wire n13643;
wire n13644;
wire n13645;
wire n13646;
wire n13647;
wire n13648;
wire n13649;
wire n13650;
wire n13651;
wire n13652;
wire n13653;
wire n13654;
wire n13655;
wire n13656;
wire n13657;
wire n13658;
wire n13659;
wire n13660;
wire n13661;
wire n13662;
wire n13663;
wire n13664;
wire n13665;
wire n13666;
wire n13667;
wire n13668;
wire n13669;
wire n13670;
wire n13671;
wire n13672;
wire n13673;
wire n13674;
wire n13675;
wire n13676;
wire n13677;
wire n13678;
wire n13679;
wire n13680;
wire n13681;
wire n13682;
wire n13683;
wire n13684;
wire n13685;
wire n13686;
wire n13687;
wire n13688;
wire n13689;
wire n13690;
wire n13691;
wire n13692;
wire n13693;
wire n13694;
wire n13695;
wire n13696;
wire n13697;
wire n13698;
wire n13699;
wire n13700;
wire n13701;
wire n13702;
wire n13703;
wire n13704;
wire n13705;
wire n13706;
wire n13707;
wire n13708;
wire n13709;
wire n13710;
wire n13711;
wire n13712;
wire n13713;
wire n13714;
wire n13715;
wire n13716;
wire n13717;
wire n13718;
wire n13719;
wire n13720;
wire n13721;
wire n13722;
wire n13723;
wire n13724;
wire n13725;
wire n13726;
wire n13727;
wire n13728;
wire n13729;
wire n13730;
wire n13731;
wire n13732;
wire n13733;
wire n13734;
wire n13735;
wire n13736;
wire n13737;
wire n13738;
wire n13739;
wire n13740;
wire n13741;
wire n13742;
wire n13743;
wire n13744;
wire n13745;
wire n13746;
wire n13747;
wire n13748;
wire n13749;
wire n13750;
wire n13751;
wire n13752;
wire n13753;
wire n13754;
wire n13755;
wire n13756;
wire n13757;
wire n13758;
wire n13759;
wire n13760;
wire n13761;
wire n13762;
wire n13763;
wire n13764;
wire n13766;
wire n13767;
wire n13768;
wire n13769;
wire n13770;
wire n13771;
wire n13772;
wire n13773;
wire n13774;
wire n13775;
wire n13776;
wire n13777;
wire n13778;
wire n13779;
wire n13780;
wire n13781;
wire n13782;
wire n13783;
wire n13784;
wire n13785;
wire n13786;
wire n13787;
wire n13788;
wire n13789;
wire n13790;
wire n13791;
wire n13792;
wire n13793;
wire n13794;
wire n13795;
wire n13796;
wire n13797;
wire n13798;
wire n13799;
wire n13800;
wire n13801;
wire n13802;
wire n13803;
wire n13804;
wire n13805;
wire n13807;
wire n13808;
wire n13809;
wire n13810;
wire n13811;
wire n13812;
wire n13813;
wire n13814;
wire n13815;
wire n13816;
wire n13817;
wire n13818;
wire n13819;
wire n13820;
wire n13821;
wire n13822;
wire n13823;
wire n13825;
wire n13826;
wire n13827;
wire n13828;
wire n13829;
wire n13830;
wire n13832;
wire n13833;
wire n13834;
wire n13835;
wire n13836;
wire n13837;
wire n13838;
wire n13839;
wire n13840;
wire n13841;
wire n13842;
wire n13843;
wire n13844;
wire n13845;
wire n13846;
wire n13847;
wire n13848;
wire n13849;
wire n13850;
wire n13853;
wire n13854;
wire n13855;
wire n13856;
wire n13857;
wire n13858;
wire n13859;
wire n13860;
wire n13861;
wire n13862;
wire n13863;
wire n13864;
wire n13865;
wire n13866;
wire n13867;
wire n13869;
wire n13870;
wire n13871;
wire n13872;
wire n13873;
wire n13874;
wire n13875;
wire n13876;
wire n13877;
wire n13878;
wire n13879;
wire n13880;
wire n13881;
wire n13882;
wire n13883;
wire n13884;
wire n13885;
wire n13886;
wire n13889;
wire n13890;
wire n13891;
wire n13894;
wire n13895;
wire n13896;
wire n13897;
wire n13898;
wire n13899;
wire n13900;
wire n13901;
wire n13903;
wire n13904;
wire n13905;
wire n13907;
wire n13908;
wire n13913;
wire n13914;
wire n13915;
wire n13916;
wire n13917;
wire n13918;
wire n13919;
wire n13920;
wire n13921;
wire NreNGPwwSfGxuZEJRmMXTmzYADEemtnb_ZN;
wire qQydNHNCopcDTmEyGIIdyrFQIErIFgJX_ZN;
wire lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN;
wire FzxTCFmmmorPYWBoKVOYVzYHHyJMkxJR_ZN;
wire rlUqTqnDczmjZLOdxrCVPPbsubqicwLv_Z;
wire KgXiNKYImGwoITNkFdnqdBmiQCHYgIoS_ZN;
wire jexoRSiRmgnTTbxiBcsGLhbKTivhVojg_Z;
wire WxUoeaFQeyYVaGStCqAbTWICyXpTFvtD_Z;

// assignments are not randomized as of now; they are copied as is
// assignments are also not considered for HD evaluation as of now, so not randomizing them does not impact the HD results

AOI21_X2 FE_RC_10_0 (.A(n11711),
.B2(n13099),
.B1(n12561),
.ZN(n12686));
INV_X8 FE_RC_9_0 (.A(FE_RN_3_0),
.ZN(n11569));
AND2_X2 FE_RC_8_0 (.A2(n11686),
.A1(n11687),
.ZN(FE_RN_3_0));
AND2_X2 FE_RC_7_0 (.A2(n11238),
.A1(n11239),
.ZN(FE_RN_2_0));
NAND3_X4 FE_RC_6_0 (.A3(n11236),
.A1(FE_RN_2_0),
.A2(n11237),
.ZN(n11428));
BUF_X1 FE_OFC32_n11469 (.A(FE_DBTN0_n11469),
.Z(FE_OFN27_n11469));
INV_X1 FE_OFC28_n11469 (.A(FE_DBTN0_n11469),
.ZN(FE_OFN23_n11469));
INV_X2 FE_OFC27_n11469 (.A(n11469),
.ZN(FE_DBTN0_n11469));
INV_X1 FE_OFC26_n12030 (.A(n12030),
.ZN(n12140));
CLKBUF_X2 FE_OFC25_n12925 (.A(n12925),
.Z(FE_OFN22_n12925));
CLKBUF_X2 FE_OFC24_n13759 (.A(n13759),
.Z(FE_OFN21_n13759));
AND2_X1 FE_RC_2_0 (.A2(n13662),
.A1(n12135),
.ZN(FE_RN_0_0));
NOR3_X1 FE_RC_1_0 (.A3(n12138),
.A1(n12888),
.A2(FE_RN_0_0),
.ZN(n12150));
XNOR2_X1 FE_RC_0_0 (.B(IR_REG_26__SCAN_IN),
.A(n11765),
.ZN(n11792));
BUF_X2 FE_OFC23_n11698 (.A(n11698),
.Z(FE_OFN20_n11698));
BUF_X1 FE_OFC19_n11466 (.A(n11466),
.Z(FE_OFN16_n11466));
INV_X2 FE_OFC18_n11466 (.A(n11466),
.ZN(n11644));
INV_X1 FE_OFC16_IR_REG_0__SCAN_IN (.A(IR_REG_0__SCAN_IN),
.ZN(n11236));
INV_X1 FE_OFC15_n11467 (.A(FE_DBTN1_n11467),
.ZN(FE_OFN14_n11467));
INV_X1 FE_OFC14_n11467 (.A(FE_DBTN1_n11467),
.ZN(FE_OFN13_n11467));
INV_X1 FE_OFC13_n11467 (.A(FE_DBTN1_n11467),
.ZN(FE_OFN12_n11467));
INV_X1 FE_OFC12_n11467 (.A(FE_DBTN1_n11467),
.ZN(FE_OFN11_n11467));
INV_X2 FE_OFC11_n11467 (.A(n11467),
.ZN(FE_DBTN1_n11467));
CLKBUF_X2 FE_OFC10_n13571 (.A(n13571),
.Z(FE_OFN10_n13571));
BUF_X1 FE_OFC9_n13503 (.A(n13503),
.Z(FE_OFN9_n13503));
CLKBUF_X2 FE_OFC8_n11821 (.A(n11821),
.Z(FE_OFN8_n11821));
CLKBUF_X3 FE_OFC7_n13835 (.A(n13835),
.Z(FE_OFN7_n13835));
BUF_X1 FE_OFC6_n13667 (.A(n13667),
.Z(FE_OFN6_n13667));
CLKBUF_X2 FE_OFC5_n12926 (.A(n12926),
.Z(FE_OFN5_n12926));
CLKBUF_X3 FE_OFC3_n13832 (.A(n13832),
.Z(FE_OFN3_n13832));
BUF_X1 FE_OFC2_n13580 (.A(n11395),
.Z(FE_OFN2_n13580));
CLKBUF_X2 FE_OFC1_n13320 (.A(n13320),
.Z(FE_OFN1_n13320));
BUF_X4 FE_OFC0_n11847 (.A(n11847),
.Z(FE_OFN0_n11847));
INV_X4 U6516 (.A(STATE_REG_SCAN_IN),
.ZN(U3149));
INV_X4 U6517 (.A(n13782),
.ZN(n11157));
INV_X1 U6521 (.A(n13138),
.ZN(n13135));
NAND2_X1 U6523 (.A2(n13189),
.A1(n13768),
.ZN(n11832));
NAND2_X1 U6524 (.A2(n13129),
.A1(n13133),
.ZN(n12434));
INV_X1 U6525 (.A(n12166),
.ZN(n12169));
INV_X1 U6527 (.A(n12423),
.ZN(n11842));
NAND2_X1 U6528 (.A2(n11336),
.A1(n11337),
.ZN(n11340));
INV_X1 U6529 (.A(n13680),
.ZN(n13214));
AND2_X1 U6531 (.A2(n11681),
.A1(n11682),
.ZN(n13768));
INV_X2 U6532 (.A(FE_OFN0_n11847),
.ZN(n11884));
NOR2_X1 U6533 (.A2(n12169),
.A1(n11832),
.ZN(n11847));
AOI21_X2 U6534 (.A(n12996),
.B2(n11908),
.B1(n12998),
.ZN(n13030));
NAND2_X1 U6535 (.A2(n11900),
.A1(n11901),
.ZN(n12998));
XNOR2_X1 U6536 (.B(n12005),
.A(n12006),
.ZN(n12120));
AOI21_X1 U6537 (.A(n11184),
.B2(n11169),
.B1(n11243),
.ZN(n11241));
NOR2_X1 U6538 (.A2(n11871),
.A1(n11872),
.ZN(n12645));
NAND2_X1 U6539 (.A2(n13123),
.A1(n13126),
.ZN(n12420));
AND2_X1 U6540 (.A2(n12429),
.A1(n11831),
.ZN(n12421));
INV_X1 U6541 (.A(n13215),
.ZN(n13700));
NAND3_X1 U6542 (.A3(n11259),
.A1(n11176),
.A2(n11377),
.ZN(n13784));
NAND2_X1 U6543 (.A2(n13315),
.A1(n13374),
.ZN(n11983));
NAND4_X1 U6544 (.A4(n11400),
.A3(n11401),
.A1(n11403),
.A2(n11402),
.ZN(n13220));
AND2_X1 U6545 (.A2(n12166),
.A1(n11832),
.ZN(n12925));
INV_X2 U6546 (.A(FE_OFN5_n12926),
.ZN(n11975));
OAI21_X1 U6547 (.A(n11368),
.B2(n11369),
.B1(n11569),
.ZN(n13128));
INV_X1 U6551 (.A(n11166),
.ZN(n12155));
AOI21_X1 U6552 (.A(n12119),
.B2(FE_OFN9_n13503),
.B1(n12120),
.ZN(n12121));
NAND2_X1 U6553 (.A2(n12004),
.A1(n12003),
.ZN(n12118));
AOI21_X1 U6554 (.A(n11693),
.B2(n13672),
.B1(n11694),
.ZN(n11807));
OAI21_X1 U6555 (.A(n12128),
.B2(n11273),
.B1(n12129),
.ZN(n12135));
OAI21_X1 U6558 (.A(n13182),
.B2(n13064),
.B1(n12006),
.ZN(n11670));
NAND2_X1 U6559 (.A2(n11261),
.A1(n11262),
.ZN(n12127));
AOI21_X1 U6560 (.A(n13356),
.B2(n13672),
.B1(n13357),
.ZN(n13601));
AOI21_X1 U6561 (.A(n12101),
.B2(n12102),
.B1(n13010),
.ZN(n12106));
AOI21_X1 U6562 (.A(n12045),
.B2(n13672),
.B1(n12046),
.ZN(n13331));
NAND2_X1 U6563 (.A2(n13062),
.A1(n11210),
.ZN(n12006));
AOI211_X1 U6565 (.C1(n13842),
.A(n13327),
.C2(n13328),
.B(n13326),
.ZN(n13329));
OAI21_X1 U6566 (.A(n12015),
.B2(FE_OFN21_n13759),
.B1(n12157),
.ZN(n12016));
AOI211_X1 U6567 (.C1(n13196),
.A(qQydNHNCopcDTmEyGIIdyrFQIErIFgJX_ZN),
.C2(n13199),
.B(n13068),
.ZN(n13194));
OAI22_X1 U6569 (.B2(n12156),
.B1(n13841),
.A1(n12157),
.A2(FE_OFN7_n13835),
.ZN(n12158));
XNOR2_X1 U6571 (.B(n13196),
.A(n12864),
.ZN(n12858));
NOR2_X1 U6573 (.A2(n13196),
.A1(n12864),
.ZN(n12866));
NAND2_X1 U6574 (.A2(n11801),
.A1(n12012),
.ZN(n12864));
NAND2_X1 U6576 (.A2(n11726),
.A1(n13479),
.ZN(n13468));
INV_X1 U6577 (.A(n12009),
.ZN(n11167));
NAND2_X1 U6578 (.A2(n11724),
.A1(n13511),
.ZN(n13480));
NOR2_X1 U6579 (.A2(n13360),
.A1(n13358),
.ZN(n11798));
NAND2_X1 U6580 (.A2(n11313),
.A1(n11723),
.ZN(n13511));
NAND2_X1 U6581 (.A2(n11661),
.A1(n11662),
.ZN(n13210));
AND2_X1 U6582 (.A2(n13395),
.A1(n13392),
.ZN(n13373));
AND2_X2 U6583 (.A2(n11193),
.A1(n13490),
.ZN(n13406));
NAND2_X1 U6584 (.A2(n11240),
.A1(n11241),
.ZN(n12614));
AND2_X1 U6585 (.A2(n13670),
.A1(n13535),
.ZN(n13490));
NAND2_X1 U6586 (.A2(n11703),
.A1(n12459),
.ZN(n11164));
AND2_X1 U6587 (.A2(n13566),
.A1(n13561),
.ZN(n13562));
AND2_X1 U6588 (.A2(n13384),
.A1(n13614),
.ZN(n11735));
OAI21_X1 U6589 (.A(n13129),
.B2(n11383),
.B1(n12435),
.ZN(n12457));
INV_X1 U6590 (.A(n11160),
.ZN(n11159));
OAI21_X1 U6591 (.A(n13486),
.B2(n11161),
.B1(n11313),
.ZN(n11160));
NAND2_X1 U6592 (.A2(n12434),
.A1(n12433),
.ZN(n11165));
NOR2_X1 U6593 (.A2(n13698),
.A1(n11157),
.ZN(n11821));
AND2_X1 U6594 (.A2(n11840),
.A1(n12263),
.ZN(n12310));
OR2_X1 U6595 (.A2(n11868),
.A1(n11869),
.ZN(n12538));
NAND2_X2 U6596 (.A2(n11993),
.A1(n13779),
.ZN(n13037));
AND2_X1 U6597 (.A2(n13094),
.A1(n11702),
.ZN(n11703));
INV_X1 U6598 (.A(n11724),
.ZN(n11161));
OAI21_X1 U6599 (.A(n12323),
.B2(n12325),
.B1(n12372),
.ZN(n12348));
NAND2_X1 U6601 (.A2(n13141),
.A1(n13136),
.ZN(n13094));
INV_X1 U6602 (.A(n13221),
.ZN(n13818));
INV_X1 U6603 (.A(n12794),
.ZN(n13216));
AND4_X1 U6606 (.A4(n11488),
.A3(n11489),
.A1(n11491),
.A2(n11490),
.ZN(n13680));
NAND2_X1 U6607 (.A2(n13215),
.A1(n12718),
.ZN(n13151));
NAND4_X1 U6608 (.A4(n11385),
.A3(n11386),
.A1(n11388),
.A2(n11387),
.ZN(n13221));
NAND2_X1 U6610 (.A2(n11314),
.A1(n11473),
.ZN(n13215));
INV_X1 U6611 (.A(n13220),
.ZN(n12618));
OR2_X1 U6612 (.A2(n12642),
.A1(FE_OFN12_n11467),
.ZN(n11423));
OR2_X1 U6613 (.A2(n12818),
.A1(n11466),
.ZN(n11478));
NAND2_X1 U6614 (.A2(n13220),
.A1(n11795),
.ZN(n13136));
INV_X1 U6615 (.A(n11260),
.ZN(n11259));
INV_X1 U6616 (.A(n12429),
.ZN(n12863));
INV_X1 U6618 (.A(n13128),
.ZN(n13132));
INV_X1 U6621 (.A(n11865),
.ZN(n12620));
INV_X1 U6624 (.A(n12822),
.ZN(n13699));
OR2_X1 U6625 (.A2(n11376),
.A1(n11418),
.ZN(n11377));
INV_X1 U6626 (.A(n13769),
.ZN(n13315));
INV_X1 U6627 (.A(n12543),
.ZN(n11795));
NAND2_X1 U6628 (.A2(n13766),
.A1(n11772),
.ZN(n12166));
INV_X1 U6630 (.A(n11792),
.ZN(n13766));
INV_X1 U6631 (.A(n13762),
.ZN(n11341));
NAND2_X1 U6633 (.A2(IR_REG_31__SCAN_IN),
.A1(n11336),
.ZN(n11332));
NOR2_X1 U6634 (.A2(IR_REG_16__SCAN_IN),
.A1(n11513),
.ZN(n11543));
NOR2_X1 U6635 (.A2(IR_REG_20__SCAN_IN),
.A1(n11671),
.ZN(n11676));
NAND2_X1 U6636 (.A2(n11177),
.A1(n11355),
.ZN(n11197));
NAND2_X1 U6637 (.A2(n11678),
.A1(IR_REG_31__SCAN_IN),
.ZN(n11679));
AND3_X1 U6638 (.A3(n11318),
.A1(n11320),
.A2(n11319),
.ZN(n11545));
NOR3_X1 U6639 (.A3(IR_REG_26__SCAN_IN),
.A1(IR_REG_28__SCAN_IN),
.A2(IR_REG_27__SCAN_IN),
.ZN(n11333));
NOR3_X1 U6640 (.A3(IR_REG_21__SCAN_IN),
.A1(IR_REG_20__SCAN_IN),
.A2(IR_REG_22__SCAN_IN),
.ZN(n11321));
INV_X1 U6641 (.A(IR_REG_7__SCAN_IN),
.ZN(n11429));
NOR2_X1 U6642 (.A2(IR_REG_5__SCAN_IN),
.A1(IR_REG_6__SCAN_IN),
.ZN(n11238));
INV_X1 U6643 (.A(IR_REG_9__SCAN_IN),
.ZN(n11451));
INV_X1 U6644 (.A(IR_REG_12__SCAN_IN),
.ZN(n11322));
INV_X1 U6645 (.A(IR_REG_11__SCAN_IN),
.ZN(n11323));
INV_X1 U6646 (.A(IR_REG_10__SCAN_IN),
.ZN(n11324));
NOR2_X1 U6648 (.A2(IR_REG_17__SCAN_IN),
.A1(IR_REG_14__SCAN_IN),
.ZN(n11320));
NOR2_X1 U6649 (.A2(IR_REG_19__SCAN_IN),
.A1(IR_REG_18__SCAN_IN),
.ZN(n11318));
NOR2_X1 U6650 (.A2(IR_REG_1__SCAN_IN),
.A1(IR_REG_2__SCAN_IN),
.ZN(n11239));
NOR2_X1 U6651 (.A2(IR_REG_15__SCAN_IN),
.A1(IR_REG_16__SCAN_IN),
.ZN(n11319));
OAI21_X2 U6652 (.A(n11159),
.B2(n11161),
.B1(n11723),
.ZN(n13479));
NAND2_X2 U6653 (.A2(n11341),
.A1(n11340),
.ZN(n11418));
NAND2_X1 U6654 (.A2(n13762),
.A1(n11340),
.ZN(n11469));
XNOR2_X1 U6655 (.B(IR_REG_30__SCAN_IN),
.A(n11332),
.ZN(n13762));
NAND3_X1 U6656 (.A3(n11256),
.A1(n11164),
.A2(n11704),
.ZN(n12506));
NAND2_X1 U6657 (.A2(n11701),
.A1(n11165),
.ZN(n12459));
NAND2_X1 U6659 (.A2(n11263),
.A1(n11737),
.ZN(n11262));
AOI21_X2 U6660 (.A(n11735),
.B2(n13376),
.B1(n13372),
.ZN(n11737));
OAI211_X1 U6661 (.C1(n12118),
.A(n12010),
.C2(n13619),
.B(n11167),
.ZN(n11166));
AOI21_X1 U6662 (.A(n12047),
.B2(n13829),
.B1(n13322),
.ZN(n12149));
XNOR2_X2 U6663 (.B(IR_REG_27__SCAN_IN),
.A(n11353),
.ZN(n11687));
NOR2_X1 U6664 (.A2(n11327),
.A1(n11673),
.ZN(n11759));
INV_X2 U6665 (.A(n11841),
.ZN(n11358));
OAI21_X2 U6666 (.A(n11364),
.B2(n11236),
.B1(n11569),
.ZN(n12429));
OAI22_X2 U6667 (.B2(n13407),
.B1(n13427),
.A1(n13416),
.A2(n11732),
.ZN(n13389));
OAI21_X1 U6668 (.A(n11832),
.B2(n11838),
.B1(n13769),
.ZN(n12926));
AND2_X1 U6669 (.A2(n13768),
.A1(n13767),
.ZN(n12168));
INV_X1 U6672 (.A(n11633),
.ZN(n11621));
NOR2_X1 U6673 (.A2(n11273),
.A1(n13117),
.ZN(n11272));
NOR2_X1 U6674 (.A2(n11613),
.A1(n11614),
.ZN(n11202));
NAND2_X1 U6677 (.A2(n12248),
.A1(n12249),
.ZN(n12251));
NAND2_X1 U6678 (.A2(REG3_REG_25__SCAN_IN),
.A1(n11202),
.ZN(n11633));
INV_X1 U6679 (.A(n11202),
.ZN(n11631));
INV_X1 U6680 (.A(n13656),
.ZN(n11915));
NOR2_X1 U6682 (.A2(n12757),
.A1(n11294),
.ZN(n11293));
NOR2_X1 U6684 (.A2(IR_REG_25__SCAN_IN),
.A1(n12197),
.ZN(n11334));
AND2_X1 U6686 (.A2(n11254),
.A1(n11448),
.ZN(n11546));
AND2_X1 U6687 (.A2(n11510),
.A1(n11255),
.ZN(n11254));
NAND2_X1 U6688 (.A2(FE_OFN5_n12926),
.A1(n11839),
.ZN(n11840));
NOR2_X1 U6689 (.A2(n12314),
.A1(n11989),
.ZN(n11997));
AOI21_X1 U6693 (.A(n11183),
.B2(n11265),
.B1(n11263),
.ZN(n11261));
AND2_X1 U6696 (.A2(n13189),
.A1(n12234),
.ZN(n13374));
INV_X2 U6697 (.A(n13690),
.ZN(n13627));
INV_X1 U6699 (.A(n12601),
.ZN(n11251));
NOR2_X1 U6700 (.A2(n12601),
.A1(n12600),
.ZN(n11252));
AOI21_X1 U6703 (.A(n12296),
.B2(n12294),
.B1(n11197),
.ZN(n12179));
NOR2_X1 U6704 (.A2(n11474),
.A1(n11475),
.ZN(n11484));
NAND2_X1 U6706 (.A2(n12309),
.A1(n12310),
.ZN(n11853));
NAND2_X1 U6707 (.A2(n12940),
.A1(n12942),
.ZN(n11250));
NOR2_X1 U6708 (.A2(n11944),
.A1(n12941),
.ZN(n11249));
NAND2_X1 U6709 (.A2(n11201),
.A1(n13225),
.ZN(n12181));
NAND2_X1 U6710 (.A2(n12774),
.A1(n12775),
.ZN(n13287));
AND2_X1 U6713 (.A2(n11640),
.A1(n11203),
.ZN(n13060));
NAND2_X1 U6714 (.A2(n13324),
.A1(n13211),
.ZN(n13059));
INV_X1 U6715 (.A(n11264),
.ZN(n11263));
OAI21_X1 U6716 (.A(n11739),
.B2(n11265),
.B1(n11736),
.ZN(n11264));
OR2_X1 U6717 (.A2(n13423),
.A1(n13089),
.ZN(n13166));
INV_X1 U6718 (.A(n13164),
.ZN(n11233));
NAND2_X1 U6719 (.A2(n11211),
.A1(n11213),
.ZN(n13048));
AOI21_X1 U6720 (.A(n11212),
.B2(n11217),
.B1(n11215),
.ZN(n11211));
INV_X1 U6721 (.A(n13156),
.ZN(n11212));
NAND2_X1 U6722 (.A2(n13154),
.A1(n13156),
.ZN(n12807));
NAND2_X1 U6723 (.A2(n12543),
.A1(n12618),
.ZN(n13141));
NAND2_X1 U6724 (.A2(n11842),
.A1(n11841),
.ZN(n13126));
NOR3_X1 U6727 (.A3(n11300),
.A1(n13335),
.A2(n11299),
.ZN(n12011));
OR2_X1 U6728 (.A2(n11974),
.A1(n12889),
.ZN(n11299));
NAND2_X1 U6729 (.A2(n13337),
.A1(n12032),
.ZN(n11300));
OR2_X1 U6730 (.A2(n13349),
.A1(n13348),
.ZN(n13377));
INV_X1 U6735 (.A(n11673),
.ZN(n11674));
AOI21_X1 U6737 (.A(n11834),
.B2(n11831),
.B1(n11846),
.ZN(n12265));
NAND2_X1 U6739 (.A2(REG3_REG_21__SCAN_IN),
.A1(n11580),
.ZN(n11601));
INV_X1 U6740 (.A(n11599),
.ZN(n11580));
NAND2_X1 U6741 (.A2(REG3_REG_15__SCAN_IN),
.A1(n11516),
.ZN(n11519));
AND2_X1 U6742 (.A2(n11632),
.A1(n11633),
.ZN(n12064));
NAND2_X1 U6743 (.A2(n11195),
.A1(n12270),
.ZN(n12283));
NAND2_X1 U6744 (.A2(n12579),
.A1(n12580),
.ZN(n12661));
AND2_X1 U6748 (.A2(n11615),
.A1(n11631),
.ZN(n13338));
INV_X1 U6750 (.A(n11229),
.ZN(n11228));
OAI21_X1 U6751 (.A(n13054),
.B2(n11230),
.B1(n11233),
.ZN(n11229));
INV_X1 U6752 (.A(n13468),
.ZN(n11279));
NAND2_X1 U6754 (.A2(n11284),
.A1(n11728),
.ZN(n11283));
INV_X1 U6755 (.A(n11727),
.ZN(n11284));
AOI21_X1 U6756 (.A(n11219),
.B2(n13150),
.B1(n11220),
.ZN(n11218));
INV_X1 U6757 (.A(n13151),
.ZN(n11219));
NAND2_X1 U6758 (.A2(n13150),
.A1(n12684),
.ZN(n11214));
INV_X1 U6759 (.A(n12807),
.ZN(n13095));
NAND2_X1 U6760 (.A2(n11714),
.A1(n11715),
.ZN(n12811));
INV_X1 U6761 (.A(n11173),
.ZN(n11220));
NAND2_X1 U6762 (.A2(REG3_REG_5__SCAN_IN),
.A1(n11397),
.ZN(n11407));
NAND2_X1 U6763 (.A2(n12429),
.A1(n12424),
.ZN(n13122));
INV_X1 U6764 (.A(n13672),
.ZN(n13568));
NAND2_X1 U6765 (.A2(n13114),
.A1(n12002),
.ZN(n12004));
NAND2_X1 U6766 (.A2(n13181),
.A1(n13065),
.ZN(n13115));
NOR2_X1 U6768 (.A2(n13586),
.A1(n13335),
.ZN(n12139));
AND2_X1 U6770 (.A2(DATAI_20_),
.A1(n11569),
.ZN(n13624));
INV_X1 U6771 (.A(n13605),
.ZN(n13628));
NAND2_X1 U6772 (.A2(n12718),
.A1(n11293),
.ZN(n11292));
INV_X1 U6773 (.A(n12677),
.ZN(n12629));
AND2_X2 U6776 (.A2(n11686),
.A1(n12168),
.ZN(n13690));
INV_X1 U6777 (.A(IR_REG_24__SCAN_IN),
.ZN(n11316));
INV_X1 U6778 (.A(IR_REG_20__SCAN_IN),
.ZN(n11683));
NAND2_X1 U6779 (.A2(IR_REG_31__SCAN_IN),
.A1(n11671),
.ZN(n11684));
NAND2_X1 U6781 (.A2(n12784),
.A1(n12785),
.ZN(n11900));
NAND2_X1 U6783 (.A2(n11245),
.A1(n11981),
.ZN(n11982));
INV_X2 U6784 (.A(n13005),
.ZN(n13043));
OR2_X1 U6786 (.A2(FE_OFN16_n11466),
.A1(n12934),
.ZN(n11662));
NAND2_X1 U6792 (.A2(n12136),
.A1(n12137),
.ZN(n12888));
INV_X1 U6793 (.A(n12134),
.ZN(n12137));
NAND2_X1 U6794 (.A2(n12452),
.A1(n12135),
.ZN(n12136));
OAI22_X1 U6795 (.B2(n12132),
.B1(n13627),
.A1(n12133),
.A2(n13568),
.ZN(n12134));
INV_X2 U6796 (.A(FE_OFN2_n13580),
.ZN(n13844));
OR2_X2 U6797 (.A2(n12314),
.A1(n11990),
.ZN(n13779));
OR2_X1 U6798 (.A2(FE_OFN7_n13835),
.A1(n12892),
.ZN(n12152));
OR2_X2 U6799 (.A2(n12027),
.A1(n12028),
.ZN(n13839));
OAI21_X1 U6800 (.A(n11268),
.B2(n11269),
.B1(n12129),
.ZN(n11267));
INV_X1 U6801 (.A(n13117),
.ZN(n11269));
NAND2_X1 U6802 (.A2(n13777),
.A1(n13226),
.ZN(n11201));
OR2_X1 U6803 (.A2(n12032),
.A1(n13212),
.ZN(n11205));
AOI21_X1 U6804 (.A(n11186),
.B2(n11216),
.B1(n11218),
.ZN(n11215));
INV_X1 U6806 (.A(n11218),
.ZN(n11217));
NAND2_X1 U6807 (.A2(n13687),
.A1(n13699),
.ZN(n13156));
NOR2_X1 U6808 (.A2(n11208),
.A1(n11561),
.ZN(n11209));
NAND2_X1 U6809 (.A2(REG3_REG_19__SCAN_IN),
.A1(REG3_REG_18__SCAN_IN),
.ZN(n11208));
NOR2_X1 U6810 (.A2(n11590),
.A1(n11601),
.ZN(n11581));
NOR2_X1 U6811 (.A2(n11506),
.A1(n11519),
.ZN(n11536));
NOR2_X1 U6812 (.A2(n11206),
.A1(n11499),
.ZN(n11516));
NAND2_X1 U6813 (.A2(REG3_REG_13__SCAN_IN),
.A1(REG3_REG_14__SCAN_IN),
.ZN(n11206));
AOI211_X1 U6814 (.C1(n13185),
.A(n13184),
.C2(n11235),
.B(n13183),
.ZN(n13186));
AOI21_X1 U6816 (.A(n12299),
.B2(n12297),
.B1(n11197),
.ZN(n12175));
NAND2_X1 U6817 (.A2(n13704),
.A1(n12571),
.ZN(n12570));
OAI21_X1 U6818 (.A(n12575),
.B2(REG1_REG_12__SCAN_IN),
.B1(n13250),
.ZN(n12577));
INV_X1 U6819 (.A(n11569),
.ZN(n12172));
INV_X1 U6820 (.A(n11738),
.ZN(n11265));
NAND2_X1 U6822 (.A2(n11713),
.A1(n13098),
.ZN(n11715));
INV_X1 U6823 (.A(n11396),
.ZN(n11397));
INV_X1 U6824 (.A(n13784),
.ZN(n11381));
NAND2_X1 U6825 (.A2(n13784),
.A1(n11382),
.ZN(n13129));
INV_X1 U6826 (.A(n13114),
.ZN(n12005));
AND2_X1 U6827 (.A2(n11298),
.A1(n13643),
.ZN(n11297));
NOR2_X1 U6828 (.A2(FzxTCFmmmorPYWBoKVOYVzYHHyJMkxJR_ZN),
.A1(n12976),
.ZN(n11298));
INV_X1 U6830 (.A(n13768),
.ZN(n13091));
INV_X1 U6831 (.A(n11209),
.ZN(n11573));
NAND2_X1 U6832 (.A2(REG3_REG_20__SCAN_IN),
.A1(n11209),
.ZN(n11599));
NAND2_X1 U6833 (.A2(REG3_REG_12__SCAN_IN),
.A1(n11484),
.ZN(n11499));
INV_X1 U6834 (.A(n11581),
.ZN(n11592));
NOR2_X1 U6836 (.A2(n11315),
.A1(n11854),
.ZN(n12386));
OR2_X1 U6837 (.A2(n11851),
.A1(n11852),
.ZN(n11854));
NAND2_X1 U6838 (.A2(REG3_REG_17__SCAN_IN),
.A1(n11536),
.ZN(n11561));
OR2_X1 U6841 (.A2(n12804),
.A1(FE_OFN14_n11467),
.ZN(n11471));
NAND2_X1 U6843 (.A2(n12463),
.A1(n12253),
.ZN(n12269));
NAND2_X1 U6844 (.A2(REG1_REG_4__SCAN_IN),
.A1(n11196),
.ZN(n12270));
OR2_X1 U6849 (.A2(n13114),
.A1(n12002),
.ZN(n12003));
NAND2_X1 U6851 (.A2(n11622),
.A1(n11633),
.ZN(n11623));
AOI21_X1 U6853 (.A(n13075),
.B2(n11225),
.B1(n11228),
.ZN(n11224));
NAND2_X1 U6854 (.A2(n11227),
.A1(n11228),
.ZN(n11226));
AND2_X1 U6855 (.A2(n11227),
.A1(n11230),
.ZN(n11225));
AOI21_X1 U6856 (.A(n11181),
.B2(n11276),
.B1(n11277),
.ZN(n11275));
INV_X1 U6857 (.A(n11175),
.ZN(n11276));
NAND2_X1 U6858 (.A2(n11233),
.A1(n11234),
.ZN(n11232));
OR2_X1 U6860 (.A2(n13547),
.A1(n13504),
.ZN(n13507));
INV_X1 U6862 (.A(n13505),
.ZN(n13547));
NAND2_X1 U6865 (.A2(REG3_REG_7__SCAN_IN),
.A1(n11420),
.ZN(n11439));
INV_X1 U6866 (.A(n11419),
.ZN(n11420));
OAI21_X1 U6868 (.A(n11378),
.B2(n12441),
.B1(FE_OFN12_n11467),
.ZN(n11260));
AND4_X1 U6869 (.A4(n11343),
.A3(n11344),
.A1(n11346),
.A2(n11345),
.ZN(n11841));
OR2_X1 U6870 (.A2(n11342),
.A1(n11418),
.ZN(n11343));
INV_X1 U6872 (.A(n11799),
.ZN(n12932));
AND2_X1 U6874 (.A2(DATAI_23_),
.A1(n11569),
.ZN(n13360));
AND2_X1 U6875 (.A2(DATAI_22_),
.A1(n11569),
.ZN(n13604));
INV_X1 U6878 (.A(n13624),
.ZN(n13407));
NAND2_X1 U6879 (.A2(n11298),
.A1(n13490),
.ZN(n13470));
INV_X1 U6880 (.A(n13036),
.ZN(n13670));
NOR2_X1 U6881 (.A2(n13534),
.A1(n13550),
.ZN(n13535));
INV_X1 U6882 (.A(n13572),
.ZN(n13692));
NOR2_X1 U6883 (.A2(n11461),
.A1(n11301),
.ZN(n12794));
INV_X1 U6884 (.A(n11293),
.ZN(n11291));
AND2_X1 U6885 (.A2(n11795),
.A1(n13135),
.ZN(n11286));
INV_X1 U6886 (.A(n13698),
.ZN(n13623));
INV_X1 U6887 (.A(n11831),
.ZN(n12424));
INV_X1 U6888 (.A(n12027),
.ZN(n11986));
NAND2_X1 U6889 (.A2(DATAI_0_),
.A1(n11569),
.ZN(n11364));
INV_X1 U6892 (.A(n12197),
.ZN(n11257));
NAND2_X1 U6893 (.A2(n13916),
.A1(IR_REG_31__SCAN_IN),
.ZN(n11350));
NAND2_X1 U6894 (.A2(n11347),
.A1(n11758),
.ZN(n11765));
NAND2_X1 U6895 (.A2(n11773),
.A1(n11675),
.ZN(n11838));
MUX2_X1 U6896 (.S(IR_REG_22__SCAN_IN),
.A(IR_REG_31__SCAN_IN),
.B(n11672),
.Z(n11675));
INV_X1 U6897 (.A(IR_REG_21__SCAN_IN),
.ZN(n11678));
NAND2_X1 U6898 (.A2(n11678),
.A1(n11676),
.ZN(n11681));
INV_X1 U6899 (.A(n11543),
.ZN(n11567));
OR2_X1 U6900 (.A2(IR_REG_10__SCAN_IN),
.A1(n11481),
.ZN(n11492));
NOR2_X1 U6901 (.A2(IR_REG_4__SCAN_IN),
.A1(IR_REG_3__SCAN_IN),
.ZN(n11237));
INV_X1 U6902 (.A(IR_REG_4__SCAN_IN),
.ZN(n11390));
OR2_X1 U6905 (.A2(n12386),
.A1(n11243),
.ZN(n11242));
INV_X1 U6906 (.A(n13037),
.ZN(n12991));
OAI21_X1 U6910 (.A(n11893),
.B2(n11304),
.B1(n12671),
.ZN(n12603));
INV_X2 U6911 (.A(n12990),
.ZN(n13038));
AOI22_X1 U6913 (.B2(n13198),
.B1(n13199),
.A1(n13201),
.A2(n13200),
.ZN(n13202));
INV_X1 U6914 (.A(n12935),
.ZN(n13211));
INV_X1 U6917 (.A(n13341),
.ZN(n13587));
INV_X1 U6918 (.A(n13614),
.ZN(n13362));
NAND2_X1 U6920 (.A2(n11554),
.A1(n11555),
.ZN(n13464));
OR2_X1 U6921 (.A2(FE_OFN16_n11466),
.A1(n13453),
.ZN(n11555));
OAI211_X1 U6922 (.C1(n13492),
.A(n11509),
.C2(FE_OFN16_n11466),
.B(n11508),
.ZN(n13667));
OR2_X1 U6925 (.A2(n11395),
.A1(n11469),
.ZN(n11401));
NOR2_X1 U6934 (.A2(n12039),
.A1(n12040),
.ZN(n12041));
AND2_X1 U6935 (.A2(n12877),
.A1(n13212),
.ZN(n12039));
INV_X1 U6937 (.A(FE_OFN8_n11821),
.ZN(n13518));
NAND2_X1 U6938 (.A2(n11231),
.A1(n13481),
.ZN(n11223));
NAND2_X1 U6941 (.A2(n11727),
.A1(n13468),
.ZN(n11280));
NAND2_X1 U6942 (.A2(n13153),
.A1(n11222),
.ZN(n12808));
NAND2_X1 U6943 (.A2(n11218),
.A1(n11214),
.ZN(n11222));
OAI21_X1 U6944 (.A(n11703),
.B2(n12477),
.B1(n12459),
.ZN(n12476));
INV_X2 U6945 (.A(n13779),
.ZN(n13842));
OR2_X1 U6946 (.A2(n11811),
.A1(n11812),
.ZN(n11809));
NOR2_X1 U6947 (.A2(n11755),
.A1(n11756),
.ZN(n11757));
NOR3_X1 U6948 (.A3(n13115),
.A1(n12004),
.A2(n13619),
.ZN(n11756));
OAI21_X1 U6950 (.A(n12051),
.B2(n13324),
.B1(n12052),
.ZN(n13325));
OR2_X1 U6953 (.A2(n12817),
.A1(n13570),
.ZN(n13760));
NOR2_X1 U6954 (.A2(n12654),
.A1(n12501),
.ZN(n12564));
NAND2_X2 U6955 (.A2(n12222),
.A1(n13204),
.ZN(n13814));
AND2_X1 U6956 (.A2(n11671),
.A1(n11547),
.ZN(n13769));
MUX2_X1 U6957 (.S(IR_REG_19__SCAN_IN),
.A(IR_REG_31__SCAN_IN),
.B(n11544),
.Z(n11547));
INV_X1 U6958 (.A(n11197),
.ZN(n13778));
AND2_X1 U6959 (.A2(n11998),
.A1(n11999),
.ZN(n12000));
NAND2_X1 U6960 (.A2(n13035),
.A1(n13210),
.ZN(n11998));
NAND2_X1 U6961 (.A2(n11270),
.A1(n11271),
.ZN(n12887));
OAI21_X1 U6962 (.A(n12159),
.B2(n13839),
.B1(n12155),
.ZN(U3546));
OR2_X1 U6963 (.A2(FE_OFN7_n13835),
.A1(n12883),
.ZN(n12033));
OR2_X1 U6965 (.A2(FE_OFN21_n13759),
.A1(n12883),
.ZN(n12037));
OR2_X1 U6966 (.A2(FE_OFN21_n13759),
.A1(n12892),
.ZN(n12143));
OR2_X1 U6967 (.A2(n12411),
.A1(n11859),
.ZN(n11169));
OAI21_X1 U6968 (.A(n11224),
.B2(n11226),
.B1(n13481),
.ZN(n13348));
NOR2_X1 U6969 (.A2(IR_REG_8__SCAN_IN),
.A1(n11494),
.ZN(n11255));
AND2_X1 U6970 (.A2(n13073),
.A1(n11182),
.ZN(n11235));
INV_X1 U6971 (.A(n13150),
.ZN(n11216));
MUX2_X1 U6972 (.S(n11569),
.A(n12252),
.B(DATAI_4_),
.Z(n13138));
AND3_X1 U6973 (.A3(n11545),
.A1(n11255),
.A2(n11510),
.ZN(n11170));
AND2_X1 U6977 (.A2(n12423),
.A1(n12863),
.ZN(n12428));
NAND2_X1 U6978 (.A2(n11236),
.A1(n11239),
.ZN(n11171));
OR2_X1 U6979 (.A2(n11918),
.A1(n11919),
.ZN(n11172));
NAND2_X1 U6980 (.A2(n11170),
.A1(n11448),
.ZN(n11671));
AOI21_X1 U6981 (.A(n11718),
.B2(n11719),
.B1(n12686),
.ZN(n13504));
NAND2_X1 U6982 (.A2(n13051),
.A1(n11232),
.ZN(n13422));
NAND2_X1 U6983 (.A2(n13216),
.A1(n12827),
.ZN(n11173));
OR2_X1 U6984 (.A2(n11549),
.A1(n11561),
.ZN(n11174));
OR2_X1 U6988 (.A2(REG3_REG_3__SCAN_IN),
.A1(n11466),
.ZN(n11176));
NAND2_X1 U6990 (.A2(n11738),
.A1(n13368),
.ZN(n13332));
NAND2_X1 U6991 (.A2(n13056),
.A1(n11612),
.ZN(n13333));
NAND2_X1 U6992 (.A2(n11228),
.A1(n11223),
.ZN(n13404));
OR2_X1 U6994 (.A2(IR_REG_1__SCAN_IN),
.A1(IR_REG_0__SCAN_IN),
.ZN(n11177));
INV_X1 U6995 (.A(n13481),
.ZN(n11234));
INV_X1 U6996 (.A(n11231),
.ZN(n11230));
NOR2_X1 U6997 (.A2(n13052),
.A1(n13166),
.ZN(n11231));
AND2_X1 U6998 (.A2(n13135),
.A1(n13221),
.ZN(n11178));
AND2_X1 U6999 (.A2(REG3_REG_6__SCAN_IN),
.A1(REG3_REG_5__SCAN_IN),
.ZN(n11179));
NOR2_X1 U7001 (.A2(n13438),
.A1(n13640),
.ZN(n11181));
OAI21_X1 U7003 (.A(n11729),
.B2(n11283),
.B1(n11730),
.ZN(n11282));
AND2_X1 U7004 (.A2(n12020),
.A1(n11205),
.ZN(n11182));
AND2_X1 U7005 (.A2(n13586),
.A1(n13213),
.ZN(n11183));
AND2_X1 U7006 (.A2(n11859),
.A1(n12411),
.ZN(n11184));
INV_X1 U7009 (.A(n11863),
.ZN(n12654));
NOR2_X1 U7011 (.A2(n11282),
.A1(n11731),
.ZN(n11277));
INV_X4 U7013 (.A(n13839),
.ZN(n13841));
NOR2_X2 U7014 (.A2(n11292),
.A1(n12501),
.ZN(n12713));
NAND2_X1 U7015 (.A2(n13658),
.A1(n13490),
.ZN(n13469));
NAND2_X1 U7016 (.A2(n11296),
.A1(n11295),
.ZN(n12563));
AND2_X1 U7017 (.A2(n13407),
.A1(n13406),
.ZN(n13392));
INV_X1 U7018 (.A(n13074),
.ZN(n11227));
OAI22_X1 U7019 (.B2(n13135),
.B1(n13221),
.A1(n12457),
.A2(n11178),
.ZN(n12474));
NAND2_X1 U7020 (.A2(n13407),
.A1(n13612),
.ZN(n13170));
XOR2_X1 U7021 (.B(n12411),
.A(n12412),
.Z(n11189));
NAND2_X1 U7022 (.A2(REG3_REG_4__SCAN_IN),
.A1(REG3_REG_3__SCAN_IN),
.ZN(n11396));
NAND2_X1 U7023 (.A2(n11255),
.A1(n11448),
.ZN(n11190));
NAND2_X1 U7024 (.A2(n11179),
.A1(n11397),
.ZN(n11419));
INV_X1 U7025 (.A(n12501),
.ZN(n11295));
AND2_X1 U7026 (.A2(n11297),
.A1(n13490),
.ZN(n13431));
AND2_X1 U7027 (.A2(REG1_REG_10__SCAN_IN),
.A1(n13772),
.ZN(n11191));
INV_X1 U7028 (.A(n13643),
.ZN(n13452));
NOR2_X1 U7029 (.A2(n11291),
.A1(n12501),
.ZN(n11192));
AND2_X1 U7030 (.A2(n13633),
.A1(n11297),
.ZN(n11193));
INV_X1 U7031 (.A(n13829),
.ZN(n13619));
NAND2_X2 U7032 (.A2(n12453),
.A1(n13488),
.ZN(n13829));
XNOR2_X1 U7033 (.B(n11683),
.A(n11684),
.ZN(n13189));
INV_X1 U7034 (.A(n13189),
.ZN(n11244));
NAND2_X1 U7035 (.A2(n13135),
.A1(n12438),
.ZN(n12461));
AND2_X1 U7037 (.A2(REG1_REG_14__SCAN_IN),
.A1(n13770),
.ZN(n11194));
INV_X1 U7038 (.A(n12889),
.ZN(n12141));
AND2_X1 U7039 (.A2(DATAI_25_),
.A1(n11569),
.ZN(n12889));
INV_X1 U7040 (.A(n13337),
.ZN(n13586));
INV_X1 U7041 (.A(IR_REG_8__SCAN_IN),
.ZN(n11447));
NAND2_X1 U7042 (.A2(n12807),
.A1(n12811),
.ZN(n12812));
OAI21_X1 U7043 (.A(n11733),
.B2(n11734),
.B1(n13389),
.ZN(n13372));
NAND2_X1 U7044 (.A2(n12796),
.A1(n13700),
.ZN(n13153));
NAND2_X1 U7045 (.A2(n12252),
.A1(n12269),
.ZN(n11195));
INV_X1 U7046 (.A(n12253),
.ZN(n11196));
MUX2_X1 U7047 (.S(n11197),
.A(n12306),
.B(n12305),
.Z(n12308));
NAND3_X1 U7048 (.A3(REG1_REG_3__SCAN_IN),
.A1(n13225),
.A2(n11201),
.ZN(n12249));
INV_X1 U7049 (.A(n12019),
.ZN(n11204));
NAND3_X1 U7050 (.A3(n11204),
.A1(n11205),
.A2(n12020),
.ZN(n11203));
NAND2_X1 U7051 (.A2(n11215),
.A1(n12684),
.ZN(n11213));
OAI21_X1 U7052 (.A(n13150),
.B2(n11220),
.B1(n12684),
.ZN(n12711));
AOI21_X2 U7053 (.A(n11404),
.B2(n13136),
.B1(n12474),
.ZN(n12523));
NAND2_X1 U7054 (.A2(n13126),
.A1(n13333),
.ZN(n12130));
NAND2_X1 U7055 (.A2(n11235),
.A1(n13333),
.ZN(n11641));
NAND2_X1 U7056 (.A2(n11169),
.A1(n12386),
.ZN(n11240));
AND2_X1 U7057 (.A2(n12387),
.A1(n12384),
.ZN(n11243));
XNOR2_X1 U7058 (.B(n11189),
.A(n11242),
.ZN(n12418));
NAND2_X2 U7059 (.A2(n11244),
.A1(n12234),
.ZN(n13698));
NOR2_X2 U7061 (.A2(n11955),
.A1(n11246),
.ZN(n13010));
AOI21_X1 U7062 (.A(n11247),
.B2(n11249),
.B1(n11250),
.ZN(n11246));
OAI22_X1 U7063 (.B2(n11251),
.B1(n11253),
.A1(n12603),
.A2(n11252),
.ZN(n12787));
NAND2_X1 U7064 (.A2(n13921),
.A1(n12787),
.ZN(n11901));
INV_X1 U7065 (.A(n12600),
.ZN(n11253));
NAND2_X1 U7066 (.A2(n11447),
.A1(n11448),
.ZN(n11495));
NAND2_X1 U7067 (.A2(n12477),
.A1(n11703),
.ZN(n11256));
NAND2_X1 U7068 (.A2(n11257),
.A1(n11258),
.ZN(n11336));
NAND2_X1 U7069 (.A2(n11759),
.A1(n11328),
.ZN(n12197));
OAI21_X1 U7070 (.A(n12026),
.B2(n12040),
.B1(n11267),
.ZN(n12035));
NAND2_X1 U7071 (.A2(n13117),
.A1(n11266),
.ZN(n11270));
NAND2_X1 U7072 (.A2(n12125),
.A1(n12129),
.ZN(n11266));
AOI21_X1 U7073 (.A(n13619),
.B2(n11273),
.B1(n13117),
.ZN(n11268));
NAND2_X1 U7074 (.A2(n11277),
.A1(n13468),
.ZN(n11274));
NAND2_X1 U7075 (.A2(n11275),
.A1(n11274),
.ZN(n13416));
NAND2_X1 U7076 (.A2(n11286),
.A1(n12438),
.ZN(n12480));
INV_X1 U7077 (.A(n12480),
.ZN(n11796));
NAND2_X1 U7078 (.A2(n11289),
.A1(n11758),
.ZN(n11353));
NAND2_X1 U7079 (.A2(n11350),
.A1(n11287),
.ZN(n11352));
NAND2_X1 U7080 (.A2(n11288),
.A1(n11758),
.ZN(n11287));
OR3_X1 U7081 (.A3(n11300),
.A1(n13335),
.A2(n12889),
.ZN(n12031));
NOR3_X1 U7082 (.A3(n12889),
.A1(n13335),
.A2(n13586),
.ZN(n12030));
NAND2_X1 U7086 (.A2(FE_OFN2_n13580),
.A1(n11803),
.ZN(n11829));
INV_X1 U7087 (.A(n12162),
.ZN(n11803));
NAND2_X1 U7088 (.A2(n12864),
.A1(n11802),
.ZN(n12162));
OAI21_X1 U7089 (.A(n12161),
.B2(FE_OFN7_n13835),
.B1(n12162),
.ZN(n12163));
AND2_X2 U7090 (.A2(n12925),
.A1(n11983),
.ZN(n11846));
NAND2_X1 U7091 (.A2(n13071),
.A1(n12127),
.ZN(n12128));
MUX2_X1 U7092 (.S(n11569),
.A(n13776),
.B(DATAI_3_),
.Z(n12490));
AOI21_X1 U7093 (.A(n11879),
.B2(n11880),
.B1(n12614),
.ZN(n12671));
NAND2_X1 U7094 (.A2(n13384),
.A1(n13373),
.ZN(n13358));
NAND2_X1 U7096 (.A2(n11356),
.A1(n11569),
.ZN(n11357));
NAND2_X1 U7097 (.A2(n11865),
.A1(n11796),
.ZN(n12501));
NAND2_X1 U7098 (.A2(n13128),
.A1(n12428),
.ZN(n12439));
NAND2_X1 U7099 (.A2(n11351),
.A1(n11352),
.ZN(n11686));
XNOR2_X1 U7100 (.B(n13069),
.A(n12866),
.ZN(n12876));
AOI21_X1 U7101 (.A(n11436),
.B2(n11437),
.B1(n12523),
.ZN(n12556));
NAND2_X2 U7102 (.A2(n13779),
.A1(n11809),
.ZN(n13782));
NOR2_X1 U7103 (.A2(n12760),
.A1(n11466),
.ZN(n11301));
INV_X1 U7106 (.A(n13633),
.ZN(n13438));
INV_X1 U7107 (.A(FE_OFN21_n13759),
.ZN(n13729));
AND3_X2 U7108 (.A3(n13203),
.A1(n11997),
.A2(n13690),
.ZN(n13035));
OR2_X1 U7109 (.A2(n12736),
.A1(n12732),
.ZN(n11304));
OR2_X1 U7110 (.A2(n11978),
.A1(n11979),
.ZN(n11305));
OR2_X1 U7111 (.A2(n12151),
.A1(n13841),
.ZN(n11306));
AND2_X1 U7113 (.A2(n12918),
.A1(n11305),
.ZN(n11309));
AND3_X1 U7117 (.A3(n13508),
.A1(n13484),
.A2(n11722),
.ZN(n11313));
INV_X1 U7118 (.A(IR_REG_31__SCAN_IN),
.ZN(n12198));
AND3_X1 U7119 (.A3(n11470),
.A1(n11472),
.A2(n11471),
.ZN(n11314));
INV_X1 U7120 (.A(n11192),
.ZN(n12712));
AND2_X1 U7121 (.A2(n11853),
.A1(n12311),
.ZN(n11315));
NAND4_X1 U7122 (.A4(n11322),
.A3(n11323),
.A1(n11451),
.A2(n11324),
.ZN(n11494));
AND2_X1 U7123 (.A2(n13076),
.A1(n13542),
.ZN(n13157));
INV_X1 U7126 (.A(REG3_REG_7__SCAN_IN),
.ZN(n11421));
NAND2_X1 U7128 (.A2(REG1_REG_9__SCAN_IN),
.A1(n12352),
.ZN(n12393));
OR2_X1 U7129 (.A2(REG2_REG_9__SCAN_IN),
.A1(n12360),
.ZN(n12398));
NAND2_X1 U7130 (.A2(n12772),
.A1(n12773),
.ZN(n12774));
INV_X1 U7131 (.A(n11516),
.ZN(n11526));
INV_X1 U7132 (.A(REG0_REG_29__SCAN_IN),
.ZN(n11804));
INV_X1 U7133 (.A(n11833),
.ZN(n11834));
INV_X1 U7134 (.A(n13777),
.ZN(n11369));
OR2_X1 U7135 (.A2(REG2_REG_12__SCAN_IN),
.A1(n12587),
.ZN(n13253));
NAND2_X1 U7136 (.A2(n13286),
.A1(n13287),
.ZN(n13290));
AND2_X1 U7140 (.A2(n13692),
.A1(n13699),
.ZN(n11797));
AND2_X1 U7141 (.A2(n11984),
.A1(n13204),
.ZN(n11789));
NAND2_X1 U7143 (.A2(n11769),
.A1(n12168),
.ZN(n13203));
NAND2_X1 U7146 (.A2(REG3_REG_28__SCAN_IN),
.A1(n13889),
.ZN(n11825));
OR2_X1 U7147 (.A2(D_REG_0__SCAN_IN),
.A1(n12222),
.ZN(n11794));
INV_X1 U7148 (.A(n13604),
.ZN(n13384));
INV_X1 U7149 (.A(n13679),
.ZN(n13554));
INV_X2 U7155 (.A(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.ZN(n13804));
NAND2_X1 U7158 (.A2(n12223),
.A1(n11794),
.ZN(n12027));
OR2_X1 U7159 (.A2(IR_REG_5__SCAN_IN),
.A1(n11393),
.ZN(n11414));
AND2_X1 U7161 (.A2(n12097),
.A1(n12098),
.ZN(n12099));
OR2_X2 U7163 (.A2(n13875),
.A1(n12182),
.ZN(n13313));
INV_X1 U7165 (.A(n11826),
.ZN(n11827));
INV_X1 U7167 (.A(n12158),
.ZN(n12159));
AND2_X1 U7169 (.A2(n12142),
.A1(n12143),
.ZN(n12144));
NAND2_X1 U7171 (.A2(n13374),
.A1(FE_OFN3_n13832),
.ZN(n13759));
INV_X1 U7174 (.A(n11838),
.ZN(n13767));
INV_X1 U7175 (.A(n12396),
.ZN(n13773));
AND2_X1 U7176 (.A2(n11414),
.A1(n11394),
.ZN(n13775));
OAI21_X1 U7177 (.A(n12148),
.B2(n13839),
.B1(n12149),
.ZN(U3545));
OAI21_X1 U7178 (.A(n12144),
.B2(n13860),
.B1(n12150),
.ZN(U3511));
NAND3_X1 U7179 (.A3(n11316),
.A1(n11447),
.A2(n11429),
.ZN(n11317));
NOR2_X1 U7180 (.A2(n11317),
.A1(n11428),
.ZN(n11328));
NAND2_X1 U7181 (.A2(n11321),
.A1(n11545),
.ZN(n11673));
INV_X1 U7182 (.A(n11494),
.ZN(n11326));
NOR2_X1 U7183 (.A2(IR_REG_23__SCAN_IN),
.A1(IR_REG_13__SCAN_IN),
.ZN(n11325));
NAND2_X1 U7184 (.A2(n11325),
.A1(n11326),
.ZN(n11327));
INV_X1 U7186 (.A(n11333),
.ZN(n11330));
NAND2_X1 U7188 (.A2(n11333),
.A1(n11334),
.ZN(n11351));
NAND2_X1 U7189 (.A2(IR_REG_31__SCAN_IN),
.A1(n11351),
.ZN(n11335));
INV_X1 U7191 (.A(n11340),
.ZN(n13763));
NAND2_X2 U7195 (.A2(n13762),
.A1(n13763),
.ZN(n11466));
NAND2_X1 U7196 (.A2(REG3_REG_1__SCAN_IN),
.A1(n11644),
.ZN(n11344));
INV_X1 U7197 (.A(REG0_REG_1__SCAN_IN),
.ZN(n11342));
NAND2_X1 U7198 (.A2(IR_REG_31__SCAN_IN),
.A1(n12197),
.ZN(n11758));
NAND2_X1 U7199 (.A2(IR_REG_25__SCAN_IN),
.A1(IR_REG_31__SCAN_IN),
.ZN(n11347));
NAND2_X1 U7201 (.A2(IR_REG_0__SCAN_IN),
.A1(IR_REG_31__SCAN_IN),
.ZN(n11354));
MUX2_X1 U7202 (.S(IR_REG_1__SCAN_IN),
.A(IR_REG_31__SCAN_IN),
.B(n11354),
.Z(n11355));
INV_X1 U7203 (.A(DATAI_1_),
.ZN(n11356));
OAI21_X2 U7204 (.A(n11357),
.B2(n13778),
.B1(n11569),
.ZN(n12423));
NAND2_X1 U7205 (.A2(n12423),
.A1(n11358),
.ZN(n13123));
INV_X1 U7206 (.A(REG2_REG_0__SCAN_IN),
.ZN(n12551));
INV_X1 U7207 (.A(REG0_REG_0__SCAN_IN),
.ZN(n11359));
NAND2_X1 U7209 (.A2(REG3_REG_0__SCAN_IN),
.A1(n11644),
.ZN(n11362));
INV_X1 U7210 (.A(REG1_REG_0__SCAN_IN),
.ZN(n11360));
OR2_X1 U7211 (.A2(n11360),
.A1(FE_OFN13_n11467),
.ZN(n11361));
NAND3_X1 U7212 (.A3(n11361),
.A1(n11363),
.A2(n11362),
.ZN(n11831));
OAI21_X1 U7213 (.A(n13126),
.B2(n13122),
.B1(n12420),
.ZN(n12446));
NAND2_X1 U7214 (.A2(IR_REG_31__SCAN_IN),
.A1(n11177),
.ZN(n11365));
MUX2_X1 U7215 (.S(IR_REG_2__SCAN_IN),
.A(IR_REG_31__SCAN_IN),
.B(n11365),
.Z(n11366));
NAND2_X1 U7216 (.A2(n11171),
.A1(n11366),
.ZN(n13777));
INV_X1 U7217 (.A(DATAI_2_),
.ZN(n11367));
NAND2_X1 U7218 (.A2(n11367),
.A1(n11569),
.ZN(n11368));
INV_X1 U7220 (.A(REG0_REG_2__SCAN_IN),
.ZN(n12703));
OR2_X1 U7221 (.A2(n12703),
.A1(n11418),
.ZN(n11372));
NOR2_X1 U7223 (.A2(FE_DBTN1_n11467),
.A1(REG1_REG_2__SCAN_IN),
.ZN(n11371));
NAND2_X1 U7224 (.A2(REG3_REG_2__SCAN_IN),
.A1(n11644),
.ZN(n11370));
NAND4_X1 U7225 (.A4(n11370),
.A3(n11371),
.A1(n11373),
.A2(n11372),
.ZN(n11698));
INV_X1 U7226 (.A(FE_OFN20_n11698),
.ZN(n13131));
OAI21_X1 U7227 (.A(n13131),
.B2(n13132),
.B1(n12446),
.ZN(n11375));
NAND2_X1 U7228 (.A2(n13132),
.A1(n12446),
.ZN(n11374));
NAND2_X1 U7229 (.A2(n11374),
.A1(n11375),
.ZN(n12435));
INV_X1 U7230 (.A(REG1_REG_3__SCAN_IN),
.ZN(n12441));
OR2_X1 U7232 (.A2(n12498),
.A1(n11469),
.ZN(n11378));
INV_X1 U7233 (.A(REG0_REG_3__SCAN_IN),
.ZN(n11376));
NAND2_X1 U7234 (.A2(IR_REG_31__SCAN_IN),
.A1(n11171),
.ZN(n11379));
MUX2_X1 U7235 (.S(IR_REG_3__SCAN_IN),
.A(IR_REG_31__SCAN_IN),
.B(n11379),
.Z(n11380));
NAND2_X1 U7237 (.A2(n12490),
.A1(n11381),
.ZN(n13133));
INV_X1 U7238 (.A(n13133),
.ZN(n11383));
INV_X1 U7239 (.A(n12490),
.ZN(n11382));
NAND2_X1 U7240 (.A2(IR_REG_31__SCAN_IN),
.A1(n11389),
.ZN(n11384));
XNOR2_X1 U7241 (.B(IR_REG_4__SCAN_IN),
.A(n11384),
.ZN(n12252));
OAI21_X1 U7242 (.A(n11396),
.B2(REG3_REG_4__SCAN_IN),
.B1(REG3_REG_3__SCAN_IN),
.ZN(n13780));
OR2_X1 U7243 (.A2(n13780),
.A1(n11466),
.ZN(n11388));
NAND2_X1 U7244 (.A2(REG1_REG_4__SCAN_IN),
.A1(FE_DBTN1_n11467),
.ZN(n11387));
INV_X1 U7245 (.A(REG2_REG_4__SCAN_IN),
.ZN(n13781));
OR2_X1 U7246 (.A2(n13781),
.A1(n11469),
.ZN(n11386));
INV_X1 U7247 (.A(REG0_REG_4__SCAN_IN),
.ZN(n12728));
OR2_X1 U7248 (.A2(n12728),
.A1(n11418),
.ZN(n11385));
NAND2_X1 U7250 (.A2(n11390),
.A1(n11391),
.ZN(n11393));
NAND2_X1 U7251 (.A2(IR_REG_31__SCAN_IN),
.A1(n11393),
.ZN(n11392));
MUX2_X1 U7252 (.S(IR_REG_5__SCAN_IN),
.A(IR_REG_31__SCAN_IN),
.B(n11392),
.Z(n11394));
MUX2_X1 U7253 (.S(n11569),
.A(n13775),
.B(DATAI_5_),
.Z(n12543));
INV_X1 U7254 (.A(REG1_REG_5__SCAN_IN),
.ZN(n13833));
OR2_X1 U7255 (.A2(n13833),
.A1(FE_OFN12_n11467),
.ZN(n11403));
INV_X1 U7256 (.A(REG0_REG_5__SCAN_IN),
.ZN(n13823));
OR2_X1 U7257 (.A2(n13823),
.A1(n11418),
.ZN(n11402));
INV_X1 U7258 (.A(REG2_REG_5__SCAN_IN),
.ZN(n11395));
INV_X1 U7259 (.A(REG3_REG_5__SCAN_IN),
.ZN(n11398));
NAND2_X1 U7260 (.A2(n11398),
.A1(n11396),
.ZN(n11399));
NAND2_X1 U7261 (.A2(n11399),
.A1(n11407),
.ZN(n12546));
OR2_X1 U7262 (.A2(n12546),
.A1(n11466),
.ZN(n11400));
INV_X1 U7263 (.A(n13141),
.ZN(n11404));
NAND2_X1 U7264 (.A2(REG2_REG_6__SCAN_IN),
.A1(FE_DBTN0_n11469),
.ZN(n11413));
INV_X1 U7265 (.A(REG0_REG_6__SCAN_IN),
.ZN(n11405));
OR2_X1 U7266 (.A2(n11405),
.A1(n11418),
.ZN(n11412));
INV_X1 U7267 (.A(REG3_REG_6__SCAN_IN),
.ZN(n11406));
NAND2_X1 U7268 (.A2(n11406),
.A1(n11407),
.ZN(n11408));
NAND2_X1 U7269 (.A2(n11408),
.A1(n11419),
.ZN(n12623));
OR2_X1 U7270 (.A2(n12623),
.A1(n11466),
.ZN(n11411));
OR2_X1 U7272 (.A2(n11409),
.A1(FE_OFN12_n11467),
.ZN(n11410));
NAND2_X1 U7274 (.A2(IR_REG_31__SCAN_IN),
.A1(n11414),
.ZN(n11415));
MUX2_X1 U7275 (.S(IR_REG_6__SCAN_IN),
.A(IR_REG_31__SCAN_IN),
.B(n11415),
.Z(n11416));
NAND2_X1 U7276 (.A2(n11428),
.A1(n11416),
.ZN(n12328));
INV_X1 U7277 (.A(DATAI_6_),
.ZN(n11417));
MUX2_X1 U7278 (.S(n11569),
.A(n12328),
.B(n11417),
.Z(n11865));
NAND2_X1 U7279 (.A2(n12620),
.A1(n12652),
.ZN(n13086));
INV_X2 U7280 (.A(n11418),
.ZN(n11645));
NAND2_X1 U7281 (.A2(REG0_REG_7__SCAN_IN),
.A1(n11645),
.ZN(n11426));
INV_X1 U7282 (.A(REG2_REG_7__SCAN_IN),
.ZN(n12375));
OR2_X1 U7283 (.A2(n12375),
.A1(n11469),
.ZN(n11425));
NAND2_X1 U7284 (.A2(n11421),
.A1(n11419),
.ZN(n11422));
NAND2_X1 U7285 (.A2(n11422),
.A1(n11439),
.ZN(n12657));
OR2_X1 U7286 (.A2(n12657),
.A1(n11466),
.ZN(n11424));
NAND2_X1 U7288 (.A2(IR_REG_31__SCAN_IN),
.A1(n11428),
.ZN(n11427));
MUX2_X1 U7289 (.S(IR_REG_7__SCAN_IN),
.A(IR_REG_31__SCAN_IN),
.B(n11427),
.Z(n11431));
INV_X1 U7290 (.A(n11428),
.ZN(n11430));
NAND2_X1 U7291 (.A2(n11429),
.A1(n11430),
.ZN(n11446));
INV_X1 U7293 (.A(DATAI_7_),
.ZN(n11432));
MUX2_X1 U7294 (.S(n11569),
.A(n12379),
.B(n11432),
.Z(n11863));
NAND2_X1 U7295 (.A2(n12654),
.A1(n12675),
.ZN(n13087));
AND2_X1 U7296 (.A2(n13087),
.A1(n13086),
.ZN(n11437));
NAND2_X1 U7297 (.A2(n13218),
.A1(n11863),
.ZN(n13143));
NAND2_X1 U7298 (.A2(n13143),
.A1(n13087),
.ZN(n12526));
NAND2_X1 U7300 (.A2(n13219),
.A1(n11865),
.ZN(n13139));
NAND2_X1 U7303 (.A2(REG2_REG_8__SCAN_IN),
.A1(FE_DBTN0_n11469),
.ZN(n11445));
INV_X1 U7304 (.A(REG0_REG_8__SCAN_IN),
.ZN(n12635));
OR2_X1 U7305 (.A2(n12635),
.A1(n11418),
.ZN(n11444));
INV_X1 U7306 (.A(REG3_REG_8__SCAN_IN),
.ZN(n11438));
NAND2_X1 U7307 (.A2(n11438),
.A1(n11439),
.ZN(n11440));
NAND2_X1 U7308 (.A2(n11440),
.A1(n11454),
.ZN(n12680));
OR2_X1 U7309 (.A2(n12680),
.A1(n11466),
.ZN(n11443));
INV_X1 U7310 (.A(REG1_REG_8__SCAN_IN),
.ZN(n11441));
OR2_X1 U7311 (.A2(n11441),
.A1(FE_OFN12_n11467),
.ZN(n11442));
NAND2_X1 U7312 (.A2(IR_REG_8__SCAN_IN),
.A1(n11446),
.ZN(n12201));
MUX2_X1 U7313 (.S(IR_REG_31__SCAN_IN),
.A(IR_REG_8__SCAN_IN),
.B(n12201),
.Z(n11449));
INV_X1 U7314 (.A(n11446),
.ZN(n11448));
MUX2_X1 U7316 (.S(n11569),
.A(n12357),
.B(DATAI_8_),
.Z(n12677));
NAND2_X1 U7317 (.A2(n12677),
.A1(n12828),
.ZN(n13148));
NAND2_X1 U7318 (.A2(n13217),
.A1(n12629),
.ZN(n13146));
NAND2_X1 U7319 (.A2(n13146),
.A1(n13148),
.ZN(n13099));
OAI21_X2 U7320 (.A(n13146),
.B2(n13099),
.B1(n12556),
.ZN(n12684));
NAND2_X1 U7321 (.A2(IR_REG_31__SCAN_IN),
.A1(n11495),
.ZN(n11450));
MUX2_X1 U7322 (.S(IR_REG_9__SCAN_IN),
.A(IR_REG_31__SCAN_IN),
.B(n11450),
.Z(n11452));
INV_X1 U7323 (.A(n11495),
.ZN(n11760));
NAND2_X1 U7324 (.A2(n11451),
.A1(n11760),
.ZN(n11481));
NAND2_X1 U7325 (.A2(n11481),
.A1(n11452),
.ZN(n12396));
MUX2_X1 U7326 (.S(n11569),
.A(n13773),
.B(DATAI_9_),
.Z(n12757));
INV_X1 U7327 (.A(n12757),
.ZN(n12827));
NAND2_X1 U7333 (.A2(REG1_REG_9__SCAN_IN),
.A1(FE_DBTN1_n11467),
.ZN(n11459));
INV_X1 U7334 (.A(REG0_REG_9__SCAN_IN),
.ZN(n12832));
OR2_X1 U7335 (.A2(n12832),
.A1(n11418),
.ZN(n11458));
NAND3_X1 U7336 (.A3(n11458),
.A1(n11460),
.A2(n11459),
.ZN(n11461));
NAND2_X1 U7337 (.A2(n12757),
.A1(n12794),
.ZN(n13150));
NAND2_X1 U7338 (.A2(IR_REG_31__SCAN_IN),
.A1(n11481),
.ZN(n11462));
XNOR2_X1 U7339 (.B(IR_REG_10__SCAN_IN),
.A(n11462),
.ZN(n13772));
MUX2_X1 U7340 (.S(n11569),
.A(n13772),
.B(DATAI_10_),
.Z(n12796));
INV_X1 U7341 (.A(n12796),
.ZN(n12718));
NAND2_X1 U7342 (.A2(REG0_REG_10__SCAN_IN),
.A1(n11645),
.ZN(n11473));
INV_X1 U7343 (.A(REG3_REG_10__SCAN_IN),
.ZN(n11463));
NAND2_X1 U7344 (.A2(n11463),
.A1(n11464),
.ZN(n11465));
NAND2_X1 U7345 (.A2(n11465),
.A1(n11475),
.ZN(n12744));
OR2_X1 U7346 (.A2(n12744),
.A1(n11466),
.ZN(n11472));
INV_X1 U7347 (.A(REG1_REG_10__SCAN_IN),
.ZN(n12804));
NAND2_X1 U7350 (.A2(REG2_REG_11__SCAN_IN),
.A1(FE_DBTN0_n11469),
.ZN(n11480));
OR2_X1 U7352 (.A2(n13704),
.A1(FE_OFN14_n11467),
.ZN(n11479));
INV_X1 U7353 (.A(REG3_REG_11__SCAN_IN),
.ZN(n11474));
INV_X1 U7354 (.A(n11484),
.ZN(n11486));
NAND2_X1 U7355 (.A2(n11474),
.A1(n11475),
.ZN(n11476));
NAND2_X1 U7356 (.A2(n11476),
.A1(n11486),
.ZN(n12818));
INV_X1 U7357 (.A(REG0_REG_11__SCAN_IN),
.ZN(n13757));
OR2_X1 U7358 (.A2(n13757),
.A1(n11418),
.ZN(n11477));
NAND2_X1 U7360 (.A2(IR_REG_31__SCAN_IN),
.A1(n11492),
.ZN(n11482));
XNOR2_X1 U7361 (.B(IR_REG_11__SCAN_IN),
.A(n11482),
.ZN(n13771));
MUX2_X1 U7362 (.S(n11569),
.A(n13771),
.B(DATAI_11_),
.Z(n12822));
NAND2_X1 U7363 (.A2(n12822),
.A1(n13578),
.ZN(n13154));
INV_X1 U7365 (.A(n13578),
.ZN(n13687));
NAND2_X1 U7366 (.A2(REG2_REG_12__SCAN_IN),
.A1(FE_DBTN0_n11469),
.ZN(n11491));
INV_X1 U7367 (.A(REG0_REG_12__SCAN_IN),
.ZN(n13753));
OR2_X1 U7368 (.A2(n13753),
.A1(n11418),
.ZN(n11490));
INV_X1 U7369 (.A(REG3_REG_12__SCAN_IN),
.ZN(n11485));
NAND2_X1 U7370 (.A2(n11485),
.A1(n11486),
.ZN(n11487));
NAND2_X1 U7371 (.A2(n11487),
.A1(n11499),
.ZN(n13573));
OR2_X1 U7372 (.A2(n13573),
.A1(n11466),
.ZN(n11489));
INV_X1 U7373 (.A(REG1_REG_12__SCAN_IN),
.ZN(n13696));
OR2_X1 U7374 (.A2(n13696),
.A1(FE_OFN14_n11467),
.ZN(n11488));
OAI21_X1 U7375 (.A(IR_REG_31__SCAN_IN),
.B2(IR_REG_11__SCAN_IN),
.B1(n11492),
.ZN(n11493));
XNOR2_X1 U7376 (.B(IR_REG_12__SCAN_IN),
.A(n11493),
.ZN(n12575));
MUX2_X1 U7377 (.S(n11569),
.A(n12575),
.B(DATAI_12_),
.Z(n13572));
NAND2_X1 U7378 (.A2(n13572),
.A1(n13680),
.ZN(n13049));
NAND2_X1 U7379 (.A2(n13049),
.A1(n13048),
.ZN(n13543));
NAND2_X1 U7380 (.A2(n13214),
.A1(n13692),
.ZN(n13542));
NAND2_X1 U7381 (.A2(IR_REG_31__SCAN_IN),
.A1(n11190),
.ZN(n11496));
INV_X1 U7382 (.A(IR_REG_13__SCAN_IN),
.ZN(n11510));
XNOR2_X1 U7383 (.B(n11510),
.A(n11496),
.ZN(n13269));
INV_X1 U7384 (.A(DATAI_13_),
.ZN(n11497));
MUX2_X1 U7385 (.S(n11569),
.A(n13269),
.B(n11497),
.Z(n13679));
INV_X1 U7386 (.A(REG3_REG_13__SCAN_IN),
.ZN(n11498));
NAND2_X1 U7389 (.A2(n13551),
.A1(n11644),
.ZN(n11504));
INV_X1 U7390 (.A(REG2_REG_13__SCAN_IN),
.ZN(n12589));
OR2_X1 U7391 (.A2(n12589),
.A1(FE_OFN23_n11469),
.ZN(n11503));
INV_X1 U7392 (.A(REG0_REG_13__SCAN_IN),
.ZN(n13749));
OR2_X1 U7393 (.A2(n13749),
.A1(n11418),
.ZN(n11502));
INV_X1 U7394 (.A(REG1_REG_13__SCAN_IN),
.ZN(n13684));
OR2_X1 U7395 (.A2(n13684),
.A1(FE_OFN14_n11467),
.ZN(n11501));
NAND2_X1 U7396 (.A2(n13689),
.A1(n13679),
.ZN(n13076));
NAND2_X1 U7397 (.A2(n13157),
.A1(n13543),
.ZN(n11505));
NAND2_X1 U7398 (.A2(n13554),
.A1(n13525),
.ZN(n13077));
NAND2_X1 U7399 (.A2(n13077),
.A1(n11505),
.ZN(n13481));
INV_X1 U7400 (.A(REG3_REG_14__SCAN_IN),
.ZN(n11524));
INV_X1 U7401 (.A(REG3_REG_16__SCAN_IN),
.ZN(n11506));
INV_X1 U7402 (.A(n11536),
.ZN(n11559));
NAND2_X1 U7403 (.A2(n11506),
.A1(n11519),
.ZN(n11507));
NAND2_X1 U7404 (.A2(n11507),
.A1(n11559),
.ZN(n13492));
AOI22_X1 U7405 (.B2(REG0_REG_16__SCAN_IN),
.B1(n11645),
.A1(FE_OFN27_n11469),
.A2(REG2_REG_16__SCAN_IN),
.ZN(n11509));
NAND2_X1 U7406 (.A2(REG1_REG_16__SCAN_IN),
.A1(FE_DBTN1_n11467),
.ZN(n11508));
NOR2_X1 U7407 (.A2(IR_REG_14__SCAN_IN),
.A1(IR_REG_15__SCAN_IN),
.ZN(n11511));
NAND2_X1 U7408 (.A2(n11511),
.A1(n11546),
.ZN(n11513));
NAND2_X1 U7409 (.A2(IR_REG_31__SCAN_IN),
.A1(n11513),
.ZN(n11512));
MUX2_X1 U7410 (.S(IR_REG_16__SCAN_IN),
.A(IR_REG_31__SCAN_IN),
.B(n11512),
.Z(n11514));
INV_X1 U7412 (.A(DATAI_16_),
.ZN(n11515));
MUX2_X1 U7413 (.S(n11569),
.A(n13288),
.B(n11515),
.Z(n13658));
OR2_X1 U7414 (.A2(n13658),
.A1(FE_OFN6_n13667),
.ZN(n13167));
INV_X1 U7415 (.A(REG3_REG_15__SCAN_IN),
.ZN(n11517));
NAND2_X1 U7416 (.A2(n11517),
.A1(n11526),
.ZN(n11518));
NAND2_X1 U7417 (.A2(n11518),
.A1(n11519),
.ZN(n13514));
OR2_X1 U7418 (.A2(FE_OFN16_n11466),
.A1(n13514),
.ZN(n11522));
AOI22_X1 U7419 (.B2(REG0_REG_15__SCAN_IN),
.B1(n11645),
.A1(FE_OFN27_n11469),
.A2(REG2_REG_15__SCAN_IN),
.ZN(n11521));
NAND2_X1 U7420 (.A2(REG1_REG_15__SCAN_IN),
.A1(FE_DBTN1_n11467),
.ZN(n11520));
INV_X1 U7421 (.A(n11546),
.ZN(n11532));
OAI21_X1 U7422 (.A(IR_REG_31__SCAN_IN),
.B2(IR_REG_14__SCAN_IN),
.B1(n11532),
.ZN(n11523));
XNOR2_X1 U7423 (.B(IR_REG_15__SCAN_IN),
.A(n11523),
.ZN(n12766));
MUX2_X1 U7424 (.S(n11569),
.A(n12766),
.B(DATAI_15_),
.Z(n13036));
NAND2_X1 U7425 (.A2(n13036),
.A1(n13526),
.ZN(n13485));
NAND2_X1 U7427 (.A2(n11524),
.A1(n11187),
.ZN(n11525));
NAND2_X1 U7429 (.A2(n11644),
.A1(n13537),
.ZN(n11531));
NAND2_X1 U7430 (.A2(REG1_REG_14__SCAN_IN),
.A1(FE_DBTN1_n11467),
.ZN(n11530));
INV_X1 U7433 (.A(REG0_REG_14__SCAN_IN),
.ZN(n13745));
OR2_X1 U7434 (.A2(n13745),
.A1(n11418),
.ZN(n11528));
NAND2_X1 U7435 (.A2(IR_REG_31__SCAN_IN),
.A1(n11532),
.ZN(n11533));
XNOR2_X1 U7436 (.B(IR_REG_14__SCAN_IN),
.A(n11533),
.ZN(n13770));
MUX2_X1 U7437 (.S(n11569),
.A(n13770),
.B(DATAI_14_),
.Z(n13534));
NAND2_X1 U7438 (.A2(n13534),
.A1(n13545),
.ZN(n13482));
INV_X1 U7441 (.A(n13534),
.ZN(n11911));
NAND2_X1 U7442 (.A2(n13666),
.A1(n11911),
.ZN(n11720));
INV_X1 U7443 (.A(n11720),
.ZN(n13483));
NAND2_X1 U7444 (.A2(n13658),
.A1(FE_OFN6_n13667),
.ZN(n11725));
NAND2_X1 U7446 (.A2(n13670),
.A1(n13655),
.ZN(n11721));
NAND2_X1 U7447 (.A2(n11721),
.A1(n11725),
.ZN(n13162));
AOI22_X1 U7448 (.B2(n13167),
.B1(n13162),
.A1(n13920),
.A2(n13483),
.ZN(n13051));
INV_X1 U7449 (.A(REG3_REG_18__SCAN_IN),
.ZN(n11549));
INV_X1 U7450 (.A(REG3_REG_19__SCAN_IN),
.ZN(n12913));
NAND2_X1 U7451 (.A2(n12913),
.A1(n11174),
.ZN(n11537));
NAND2_X1 U7452 (.A2(n11537),
.A1(n11573),
.ZN(n13434));
INV_X1 U7453 (.A(REG1_REG_19__SCAN_IN),
.ZN(n13638));
NAND2_X1 U7454 (.A2(REG0_REG_19__SCAN_IN),
.A1(n11645),
.ZN(n11539));
NAND2_X1 U7455 (.A2(REG2_REG_19__SCAN_IN),
.A1(FE_OFN27_n11469),
.ZN(n11538));
OAI211_X1 U7456 (.C1(FE_OFN11_n11467),
.A(n11539),
.C2(n13638),
.B(n11538),
.ZN(n11540));
INV_X1 U7457 (.A(n11540),
.ZN(n11541));
OAI21_X2 U7458 (.A(n11541),
.B2(FE_OFN16_n11466),
.B1(n13434),
.ZN(n13640));
NOR2_X1 U7459 (.A2(IR_REG_17__SCAN_IN),
.A1(IR_REG_18__SCAN_IN),
.ZN(n11542));
NAND2_X1 U7460 (.A2(n11542),
.A1(n11543),
.ZN(n12212));
NAND2_X1 U7461 (.A2(IR_REG_31__SCAN_IN),
.A1(n12212),
.ZN(n11544));
INV_X1 U7462 (.A(DATAI_19_),
.ZN(n11548));
MUX2_X1 U7463 (.S(n11569),
.A(n13315),
.B(n11548),
.Z(n13633));
NAND2_X1 U7464 (.A2(n13633),
.A1(n13640),
.ZN(n13420));
NAND2_X1 U7465 (.A2(n11549),
.A1(n11561),
.ZN(n11550));
NAND2_X1 U7466 (.A2(n11550),
.A1(n11174),
.ZN(n13453));
INV_X1 U7467 (.A(REG2_REG_18__SCAN_IN),
.ZN(n13454));
NAND2_X1 U7468 (.A2(REG1_REG_18__SCAN_IN),
.A1(FE_DBTN1_n11467),
.ZN(n11552));
NAND2_X1 U7469 (.A2(REG0_REG_18__SCAN_IN),
.A1(n11645),
.ZN(n11551));
OAI211_X1 U7470 (.C1(FE_OFN23_n11469),
.A(n11552),
.C2(n13454),
.B(n11551),
.ZN(n11553));
INV_X1 U7471 (.A(n11553),
.ZN(n11554));
OAI21_X1 U7472 (.A(IR_REG_18__SCAN_IN),
.B2(IR_REG_17__SCAN_IN),
.B1(n11567),
.ZN(n12213));
MUX2_X1 U7473 (.S(IR_REG_31__SCAN_IN),
.A(IR_REG_18__SCAN_IN),
.B(n12213),
.Z(n11556));
INV_X1 U7475 (.A(DATAI_18_),
.ZN(n11557));
MUX2_X1 U7476 (.S(n11569),
.A(n13307),
.B(n11557),
.Z(n13643));
NAND2_X1 U7477 (.A2(n13643),
.A1(n13464),
.ZN(n13443));
NAND2_X1 U7478 (.A2(n13443),
.A1(n13420),
.ZN(n13089));
INV_X1 U7479 (.A(REG3_REG_17__SCAN_IN),
.ZN(n11558));
NAND2_X1 U7480 (.A2(n11558),
.A1(n11559),
.ZN(n11560));
NAND2_X1 U7481 (.A2(n11560),
.A1(n11561),
.ZN(n13473));
NAND2_X1 U7483 (.A2(REG2_REG_17__SCAN_IN),
.A1(FE_OFN27_n11469),
.ZN(n11563));
NAND2_X1 U7484 (.A2(REG0_REG_17__SCAN_IN),
.A1(n11645),
.ZN(n11562));
OAI211_X1 U7485 (.C1(n13653),
.A(n11563),
.C2(FE_OFN11_n11467),
.B(n11562),
.ZN(n11564));
NAND2_X1 U7487 (.A2(IR_REG_31__SCAN_IN),
.A1(n11567),
.ZN(n11568));
XNOR2_X1 U7488 (.B(IR_REG_17__SCAN_IN),
.A(n11568),
.ZN(n13810));
MUX2_X1 U7489 (.S(n11569),
.A(n13810),
.B(DATAI_17_),
.Z(n12976));
INV_X1 U7490 (.A(n12976),
.ZN(n13471));
NOR2_X1 U7492 (.A2(n13643),
.A1(n13464),
.ZN(n13445));
OR2_X1 U7497 (.A2(n13424),
.A1(n13089),
.ZN(n11571));
AND2_X1 U7498 (.A2(n11571),
.A1(n11572),
.ZN(n13054));
INV_X1 U7499 (.A(REG3_REG_20__SCAN_IN),
.ZN(n12989));
NAND2_X1 U7500 (.A2(n12989),
.A1(n11573),
.ZN(n11574));
AND2_X1 U7501 (.A2(n11574),
.A1(n11599),
.ZN(n13409));
INV_X1 U7503 (.A(REG1_REG_20__SCAN_IN),
.ZN(n13631));
NAND2_X1 U7504 (.A2(REG2_REG_20__SCAN_IN),
.A1(FE_OFN27_n11469),
.ZN(n11576));
NAND2_X1 U7505 (.A2(REG0_REG_20__SCAN_IN),
.A1(n11645),
.ZN(n11575));
OAI211_X1 U7506 (.C1(n13631),
.A(n11576),
.C2(FE_OFN11_n11467),
.B(n11575),
.ZN(n11577));
NOR2_X1 U7508 (.A2(n13407),
.A1(n13612),
.ZN(n13074));
INV_X1 U7509 (.A(REG3_REG_22__SCAN_IN),
.ZN(n11590));
NAND2_X1 U7510 (.A2(REG3_REG_23__SCAN_IN),
.A1(n11581),
.ZN(n11614));
INV_X1 U7511 (.A(REG3_REG_23__SCAN_IN),
.ZN(n11582));
NAND2_X1 U7512 (.A2(n11582),
.A1(n11592),
.ZN(n11583));
NAND2_X1 U7513 (.A2(n11583),
.A1(n11614),
.ZN(n12079));
INV_X1 U7514 (.A(REG1_REG_23__SCAN_IN),
.ZN(n11586));
NAND2_X1 U7515 (.A2(REG0_REG_23__SCAN_IN),
.A1(n11645),
.ZN(n11585));
NAND2_X1 U7516 (.A2(REG2_REG_23__SCAN_IN),
.A1(FE_OFN27_n11469),
.ZN(n11584));
OAI211_X1 U7517 (.C1(FE_OFN11_n11467),
.A(n11585),
.C2(n11586),
.B(n11584),
.ZN(n11587));
NAND2_X1 U7519 (.A2(n13360),
.A1(n13341),
.ZN(n13121));
NAND2_X1 U7520 (.A2(n11590),
.A1(n11601),
.ZN(n11591));
AND2_X1 U7521 (.A2(n11591),
.A1(n11592),
.ZN(n13381));
INV_X1 U7523 (.A(REG1_REG_22__SCAN_IN),
.ZN(n11595));
NAND2_X1 U7524 (.A2(REG0_REG_22__SCAN_IN),
.A1(n11645),
.ZN(n11594));
NAND2_X1 U7525 (.A2(REG2_REG_22__SCAN_IN),
.A1(FE_OFN27_n11469),
.ZN(n11593));
OAI211_X1 U7526 (.C1(FE_OFN11_n11467),
.A(n11594),
.C2(n11595),
.B(n11593),
.ZN(n11596));
NAND2_X1 U7528 (.A2(n13604),
.A1(n13614),
.ZN(n13353));
NAND2_X1 U7529 (.A2(n13353),
.A1(n13121),
.ZN(n11608));
INV_X1 U7530 (.A(REG3_REG_21__SCAN_IN),
.ZN(n12948));
NAND2_X1 U7531 (.A2(n12948),
.A1(n11599),
.ZN(n11600));
NAND2_X1 U7532 (.A2(n11600),
.A1(n11601),
.ZN(n13398));
INV_X1 U7533 (.A(REG1_REG_21__SCAN_IN),
.ZN(n11604));
NAND2_X1 U7534 (.A2(REG2_REG_21__SCAN_IN),
.A1(FE_OFN27_n11469),
.ZN(n11603));
NAND2_X1 U7535 (.A2(REG0_REG_21__SCAN_IN),
.A1(n11645),
.ZN(n11602));
OAI211_X1 U7536 (.C1(n11604),
.A(n11603),
.C2(FE_OFN11_n11467),
.B(n11602),
.ZN(n11605));
NOR2_X1 U7538 (.A2(n13350),
.A1(n11608),
.ZN(n13173));
NAND2_X1 U7539 (.A2(n13173),
.A1(n13348),
.ZN(n11612));
INV_X1 U7540 (.A(n11608),
.ZN(n11611));
NAND2_X1 U7541 (.A2(n13384),
.A1(n13362),
.ZN(n13177));
NAND2_X1 U7542 (.A2(n13395),
.A1(n13605),
.ZN(n13169));
NAND2_X1 U7543 (.A2(n13169),
.A1(n13177),
.ZN(n11610));
INV_X1 U7544 (.A(n13360),
.ZN(n13595));
NAND2_X1 U7545 (.A2(n13595),
.A1(n13587),
.ZN(n13175));
INV_X1 U7546 (.A(n13175),
.ZN(n11609));
AOI21_X1 U7547 (.A(n11609),
.B2(n11610),
.B1(n11611),
.ZN(n13056));
INV_X1 U7548 (.A(REG3_REG_24__SCAN_IN),
.ZN(n11613));
NAND2_X1 U7549 (.A2(n11613),
.A1(n11614),
.ZN(n11615));
NAND2_X1 U7550 (.A2(n11644),
.A1(n13338),
.ZN(n11620));
INV_X1 U7551 (.A(REG1_REG_24__SCAN_IN),
.ZN(n13593));
NAND2_X1 U7552 (.A2(REG2_REG_24__SCAN_IN),
.A1(FE_OFN27_n11469),
.ZN(n11617));
NAND2_X1 U7553 (.A2(REG0_REG_24__SCAN_IN),
.A1(n11645),
.ZN(n11616));
OAI211_X1 U7554 (.C1(n13593),
.A(n11617),
.C2(FE_OFN11_n11467),
.B(n11616),
.ZN(n11618));
INV_X1 U7555 (.A(n11618),
.ZN(n11619));
NAND2_X1 U7556 (.A2(DATAI_24_),
.A1(n11569),
.ZN(n13337));
NAND2_X1 U7557 (.A2(n13586),
.A1(n13355),
.ZN(n13073));
INV_X1 U7558 (.A(REG3_REG_25__SCAN_IN),
.ZN(n11630));
NAND2_X1 U7559 (.A2(REG3_REG_26__SCAN_IN),
.A1(n11621),
.ZN(n11642));
INV_X1 U7560 (.A(REG3_REG_26__SCAN_IN),
.ZN(n11622));
NAND2_X1 U7561 (.A2(n11623),
.A1(n11642),
.ZN(n12880));
INV_X1 U7562 (.A(REG1_REG_26__SCAN_IN),
.ZN(n11626));
NAND2_X1 U7563 (.A2(REG2_REG_26__SCAN_IN),
.A1(FE_DBTN0_n11469),
.ZN(n11625));
NAND2_X1 U7564 (.A2(REG0_REG_26__SCAN_IN),
.A1(n11645),
.ZN(n11624));
OAI211_X1 U7565 (.C1(n11626),
.A(n11625),
.C2(FE_OFN11_n11467),
.B(n11624),
.ZN(n11627));
NAND2_X1 U7567 (.A2(n11630),
.A1(n11631),
.ZN(n11632));
INV_X1 U7568 (.A(REG1_REG_25__SCAN_IN),
.ZN(n12151));
NAND2_X1 U7569 (.A2(REG2_REG_25__SCAN_IN),
.A1(FE_OFN27_n11469),
.ZN(n11635));
NAND2_X1 U7570 (.A2(REG0_REG_25__SCAN_IN),
.A1(n11645),
.ZN(n11634));
OAI211_X1 U7571 (.C1(n12151),
.A(n11635),
.C2(FE_OFN11_n11467),
.B(n11634),
.ZN(n11636));
NAND2_X1 U7573 (.A2(n12889),
.A1(n13890),
.ZN(n12020));
NAND2_X1 U7577 (.A2(n12032),
.A1(n13212),
.ZN(n11640));
INV_X1 U7579 (.A(REG3_REG_27__SCAN_IN),
.ZN(n11994));
INV_X1 U7582 (.A(REG1_REG_27__SCAN_IN),
.ZN(n12145));
NAND2_X1 U7583 (.A2(REG2_REG_27__SCAN_IN),
.A1(FE_OFN27_n11469),
.ZN(n11647));
NAND2_X1 U7584 (.A2(REG0_REG_27__SCAN_IN),
.A1(n11645),
.ZN(n11646));
OAI211_X1 U7585 (.C1(FE_OFN11_n11467),
.A(n11647),
.C2(n12145),
.B(n11646),
.ZN(n11648));
NAND2_X1 U7588 (.A2(n11974),
.A1(n12935),
.ZN(n13062));
INV_X1 U7590 (.A(REG3_REG_28__SCAN_IN),
.ZN(n11653));
NAND2_X1 U7591 (.A2(n11653),
.A1(n11654),
.ZN(n11655));
NAND2_X1 U7592 (.A2(n11655),
.A1(n11825),
.ZN(n12934));
INV_X1 U7593 (.A(REG1_REG_28__SCAN_IN),
.ZN(n12156));
NAND2_X1 U7594 (.A2(REG0_REG_28__SCAN_IN),
.A1(n11645),
.ZN(n11658));
NAND2_X1 U7595 (.A2(REG2_REG_28__SCAN_IN),
.A1(FE_DBTN0_n11469),
.ZN(n11657));
OAI211_X1 U7596 (.C1(FE_OFN11_n11467),
.A(n11658),
.C2(n12156),
.B(n11657),
.ZN(n11660));
INV_X1 U7597 (.A(n11660),
.ZN(n11661));
NAND2_X1 U7598 (.A2(DATAI_28_),
.A1(n11569),
.ZN(n11799));
NOR2_X1 U7599 (.A2(n11799),
.A1(n13210),
.ZN(n13064));
NAND2_X1 U7600 (.A2(n11799),
.A1(n13210),
.ZN(n13182));
INV_X1 U7601 (.A(REG2_REG_29__SCAN_IN),
.ZN(n11666));
NAND2_X1 U7602 (.A2(REG1_REG_29__SCAN_IN),
.A1(FE_DBTN1_n11467),
.ZN(n11665));
OR2_X1 U7603 (.A2(n11804),
.A1(n11418),
.ZN(n11664));
OAI211_X1 U7604 (.C1(n11469),
.A(n11665),
.C2(n11666),
.B(n11664),
.ZN(n11667));
NAND2_X1 U7606 (.A2(DATAI_29_),
.A1(n11569),
.ZN(n11801));
NAND2_X1 U7607 (.A2(n11801),
.A1(n13209),
.ZN(n13181));
XNOR2_X1 U7608 (.B(n13115),
.A(n11670),
.ZN(n11694));
NAND2_X1 U7609 (.A2(IR_REG_31__SCAN_IN),
.A1(n11681),
.ZN(n11672));
NAND2_X1 U7610 (.A2(n11674),
.A1(n11546),
.ZN(n11773));
NAND2_X1 U7611 (.A2(n13767),
.A1(n13769),
.ZN(n11685));
NAND2_X1 U7614 (.A2(n11679),
.A1(n11680),
.ZN(n11682));
NAND2_X1 U7615 (.A2(n11244),
.A1(n13768),
.ZN(n13193));
NAND2_X1 U7618 (.A2(n11689),
.A1(n13690),
.ZN(n12843));
NAND2_X1 U7619 (.A2(REG1_REG_30__SCAN_IN),
.A1(FE_DBTN1_n11467),
.ZN(n11692));
INV_X1 U7620 (.A(REG2_REG_30__SCAN_IN),
.ZN(n12852));
OR2_X1 U7621 (.A2(n12852),
.A1(n11469),
.ZN(n11691));
INV_X1 U7622 (.A(REG0_REG_30__SCAN_IN),
.ZN(n12849));
OR2_X1 U7623 (.A2(n12849),
.A1(n11418),
.ZN(n11690));
AND3_X1 U7624 (.A3(n11690),
.A1(n11692),
.A2(n11691),
.ZN(n13197));
NOR2_X1 U7625 (.A2(n13197),
.A1(n12843),
.ZN(n11693));
NAND2_X1 U7626 (.A2(n12423),
.A1(n11841),
.ZN(n11695));
NAND2_X1 U7627 (.A2(n11695),
.A1(n12421),
.ZN(n11697));
OR2_X1 U7628 (.A2(n11841),
.A1(n12423),
.ZN(n11696));
XNOR2_X1 U7630 (.B(n13128),
.A(FE_OFN20_n11698),
.ZN(n13083));
NAND2_X1 U7631 (.A2(n13083),
.A1(n12444),
.ZN(n11700));
NAND2_X1 U7632 (.A2(FE_OFN20_n11698),
.A1(n13132),
.ZN(n11699));
NAND2_X1 U7633 (.A2(n11699),
.A1(n11700),
.ZN(n12433));
NAND2_X1 U7634 (.A2(n13784),
.A1(n12490),
.ZN(n11701));
AND2_X1 U7635 (.A2(n13221),
.A1(n13138),
.ZN(n12477));
NAND2_X1 U7636 (.A2(n13135),
.A1(n13818),
.ZN(n11702));
NAND2_X1 U7637 (.A2(n13220),
.A1(n12543),
.ZN(n11704));
AOI22_X1 U7638 (.B2(n11863),
.B1(n12675),
.A1(n12652),
.A2(n11865),
.ZN(n11705));
NAND2_X1 U7639 (.A2(n11705),
.A1(n12506),
.ZN(n11710));
NAND2_X1 U7640 (.A2(n13219),
.A1(n12620),
.ZN(n11706));
NAND2_X1 U7641 (.A2(n12675),
.A1(n11706),
.ZN(n11708));
AND2_X1 U7642 (.A2(n13218),
.A1(n13219),
.ZN(n11707));
AOI22_X1 U7643 (.B2(n12620),
.B1(n11707),
.A1(n11708),
.A2(n12654),
.ZN(n11709));
AND2_X1 U7645 (.A2(n13217),
.A1(n12677),
.ZN(n11711));
NAND2_X1 U7647 (.A2(n13216),
.A1(n12757),
.ZN(n12707));
AND2_X1 U7648 (.A2(n13153),
.A1(n13151),
.ZN(n13098));
NAND2_X1 U7649 (.A2(n12718),
.A1(n13700),
.ZN(n11713));
AND2_X1 U7650 (.A2(n11715),
.A1(n12707),
.ZN(n12810));
NAND2_X1 U7651 (.A2(n13687),
.A1(n12822),
.ZN(n11716));
AND2_X1 U7652 (.A2(n11716),
.A1(n12810),
.ZN(n13559));
NAND2_X1 U7653 (.A2(n13214),
.A1(n13572),
.ZN(n11712));
AND2_X1 U7654 (.A2(n11712),
.A1(n13559),
.ZN(n11719));
NAND2_X1 U7656 (.A2(n12794),
.A1(n12827),
.ZN(n12708));
NAND2_X1 U7657 (.A2(n11713),
.A1(n12708),
.ZN(n11714));
NAND2_X1 U7658 (.A2(n11716),
.A1(n12812),
.ZN(n13561));
NAND2_X1 U7659 (.A2(n13542),
.A1(n13049),
.ZN(n13566));
NOR2_X1 U7660 (.A2(n13562),
.A1(n11712),
.ZN(n11718));
NAND2_X1 U7661 (.A2(n11720),
.A1(n13482),
.ZN(n13524));
NAND2_X1 U7662 (.A2(n13679),
.A1(n13525),
.ZN(n13506));
NAND3_X1 U7663 (.A3(n13506),
.A1(n13504),
.A2(n13524),
.ZN(n11723));
NAND2_X1 U7664 (.A2(n11721),
.A1(n13485),
.ZN(n13484));
NAND3_X1 U7665 (.A3(n13689),
.A1(n13524),
.A2(n13554),
.ZN(n11722));
NAND2_X1 U7666 (.A2(n13666),
.A1(n13534),
.ZN(n13508));
NAND2_X1 U7667 (.A2(n13670),
.A1(n13526),
.ZN(n11724));
NAND2_X1 U7668 (.A2(n11725),
.A1(n13167),
.ZN(n13486));
INV_X1 U7669 (.A(n13658),
.ZN(n13491));
OR2_X1 U7670 (.A2(FzxTCFmmmorPYWBoKVOYVzYHHyJMkxJR_ZN),
.A1(FE_OFN6_n13667),
.ZN(n11726));
NAND2_X1 U7671 (.A2(n12976),
.A1(n13656),
.ZN(n11727));
NAND2_X1 U7672 (.A2(n13471),
.A1(n11915),
.ZN(n11728));
NOR2_X1 U7673 (.A2(n13452),
.A1(n13464),
.ZN(n11730));
NAND2_X1 U7674 (.A2(n13452),
.A1(n13464),
.ZN(n11729));
AND2_X1 U7675 (.A2(n13438),
.A1(n13640),
.ZN(n11731));
NOR2_X1 U7676 (.A2(n13624),
.A1(n13612),
.ZN(n11732));
AND2_X1 U7678 (.A2(n13611),
.A1(n13605),
.ZN(n11734));
NAND2_X1 U7679 (.A2(n13395),
.A1(n13628),
.ZN(n11733));
NAND2_X1 U7680 (.A2(n13177),
.A1(n13353),
.ZN(n13376));
NAND2_X1 U7681 (.A2(n13360),
.A1(n13587),
.ZN(n11738));
NAND2_X1 U7682 (.A2(n13337),
.A1(n13355),
.ZN(n11739));
OAI21_X1 U7683 (.A(n12125),
.B2(n12877),
.B1(n13212),
.ZN(n11740));
INV_X1 U7684 (.A(n11740),
.ZN(n11741));
NAND2_X1 U7685 (.A2(n11741),
.A1(n12127),
.ZN(n11746));
NAND2_X1 U7686 (.A2(n13059),
.A1(n13062),
.ZN(n13113));
NAND3_X1 U7687 (.A3(n12889),
.A1(n13343),
.A2(n12877),
.ZN(n11743));
OAI21_X1 U7688 (.A(n13212),
.B2(n12877),
.B1(n12124),
.ZN(n11742));
AND3_X1 U7689 (.A3(n11742),
.A1(n13113),
.A2(n11743),
.ZN(n11745));
AND2_X1 U7690 (.A2(n13324),
.A1(n12935),
.ZN(n11744));
INV_X1 U7692 (.A(n13064),
.ZN(n11747));
NAND2_X1 U7693 (.A2(n13182),
.A1(n11747),
.ZN(n13114));
INV_X1 U7694 (.A(n12168),
.ZN(n11981));
NAND2_X1 U7695 (.A2(n11838),
.A1(n11832),
.ZN(n11748));
NAND3_X1 U7696 (.A3(n11748),
.A1(n11981),
.A2(n13315),
.ZN(n13488));
NAND2_X1 U7698 (.A2(n12932),
.A1(n13210),
.ZN(n11815));
NAND4_X1 U7699 (.A4(n11815),
.A3(n13115),
.A1(n12004),
.A2(n13829),
.ZN(n11754));
NAND3_X1 U7700 (.A3(n13829),
.A1(n13210),
.A2(n12932),
.ZN(n11751));
INV_X1 U7701 (.A(n11686),
.ZN(n13764));
NOR2_X1 U7702 (.A2(n11801),
.A1(n13698),
.ZN(n11749));
AOI21_X1 U7703 (.A(n11749),
.B2(n13688),
.B1(n13210),
.ZN(n11750));
OAI21_X1 U7704 (.A(n11750),
.B2(n11751),
.B1(n13115),
.ZN(n11752));
INV_X1 U7705 (.A(n11752),
.ZN(n11753));
NAND2_X1 U7706 (.A2(n11753),
.A1(n11754),
.ZN(n11755));
NAND2_X1 U7707 (.A2(n11757),
.A1(n11807),
.ZN(n12160));
NAND2_X1 U7708 (.A2(n13091),
.A1(n13662),
.ZN(n11990));
XNOR2_X1 U7709 (.B(n11329),
.A(n11758),
.ZN(n11770));
NAND2_X1 U7710 (.A2(B_REG_SCAN_IN),
.A1(n11770),
.ZN(n11764));
NAND2_X1 U7711 (.A2(n11759),
.A1(n11760),
.ZN(n11775));
NAND2_X1 U7712 (.A2(IR_REG_24__SCAN_IN),
.A1(n11775),
.ZN(n12196));
INV_X1 U7713 (.A(n11758),
.ZN(n11761));
MUX2_X1 U7717 (.S(n11791),
.A(n11764),
.B(B_REG_SCAN_IN),
.Z(n11767));
OR2_X1 U7720 (.A2(D_REG_1__SCAN_IN),
.A1(n12222),
.ZN(n11768));
NAND2_X1 U7721 (.A2(n11770),
.A1(n11792),
.ZN(n13761));
NAND2_X1 U7722 (.A2(n13761),
.A1(n11768),
.ZN(n11808));
NAND2_X1 U7724 (.A2(n13189),
.A1(n13315),
.ZN(n11769));
NAND2_X1 U7727 (.A2(IR_REG_31__SCAN_IN),
.A1(n11773),
.ZN(n11774));
MUX2_X1 U7728 (.S(IR_REG_23__SCAN_IN),
.A(IR_REG_31__SCAN_IN),
.B(n11774),
.Z(n11776));
NOR4_X1 U7730 (.A4(D_REG_21__SCAN_IN),
.A3(D_REG_20__SCAN_IN),
.A1(D_REG_18__SCAN_IN),
.A2(D_REG_19__SCAN_IN),
.ZN(n11781));
NOR4_X1 U7731 (.A4(D_REG_17__SCAN_IN),
.A3(D_REG_15__SCAN_IN),
.A1(D_REG_16__SCAN_IN),
.A2(D_REG_14__SCAN_IN),
.ZN(n11780));
NOR4_X1 U7732 (.A4(D_REG_31__SCAN_IN),
.A3(D_REG_28__SCAN_IN),
.A1(D_REG_26__SCAN_IN),
.A2(D_REG_27__SCAN_IN),
.ZN(n11779));
NOR4_X1 U7733 (.A4(D_REG_25__SCAN_IN),
.A3(D_REG_24__SCAN_IN),
.A1(D_REG_22__SCAN_IN),
.A2(D_REG_23__SCAN_IN),
.ZN(n11778));
NAND4_X1 U7734 (.A4(n11778),
.A3(n11779),
.A1(n11781),
.A2(n11780),
.ZN(n11787));
NOR2_X1 U7735 (.A2(D_REG_3__SCAN_IN),
.A1(D_REG_2__SCAN_IN),
.ZN(n11785));
NOR4_X1 U7736 (.A4(D_REG_5__SCAN_IN),
.A3(D_REG_4__SCAN_IN),
.A1(D_REG_29__SCAN_IN),
.A2(D_REG_30__SCAN_IN),
.ZN(n11784));
NOR4_X1 U7737 (.A4(D_REG_13__SCAN_IN),
.A3(D_REG_12__SCAN_IN),
.A1(D_REG_10__SCAN_IN),
.A2(D_REG_11__SCAN_IN),
.ZN(n11783));
NOR4_X1 U7738 (.A4(D_REG_9__SCAN_IN),
.A3(D_REG_8__SCAN_IN),
.A1(D_REG_6__SCAN_IN),
.A2(D_REG_7__SCAN_IN),
.ZN(n11782));
NAND4_X1 U7739 (.A4(n11782),
.A3(n11783),
.A1(n11785),
.A2(n11784),
.ZN(n11786));
NAND2_X1 U7742 (.A2(n11792),
.A1(n13907),
.ZN(n12223));
NAND2_X1 U7744 (.A2(FE_OFN3_n13832),
.A1(n12160),
.ZN(n11806));
NAND2_X1 U7745 (.A2(n11797),
.A1(n12713),
.ZN(n13548));
OR2_X1 U7746 (.A2(n13554),
.A1(n13548),
.ZN(n13550));
INV_X1 U7747 (.A(n11798),
.ZN(n13335));
INV_X1 U7749 (.A(n11801),
.ZN(n11822));
NAND2_X1 U7750 (.A2(n11822),
.A1(n11800),
.ZN(n11802));
NAND2_X1 U7752 (.A2(n11308),
.A1(n11806),
.ZN(U3515));
INV_X1 U7753 (.A(n11807),
.ZN(n11810));
INV_X1 U7754 (.A(n11808),
.ZN(n11985));
NAND2_X1 U7755 (.A2(n12027),
.A1(n11985),
.ZN(n11811));
NAND2_X1 U7756 (.A2(n13782),
.A1(n11810),
.ZN(n11830));
NAND2_X1 U7759 (.A2(n11815),
.A1(n12004),
.ZN(n11816));
INV_X1 U7761 (.A(n11832),
.ZN(n11817));
AND2_X1 U7762 (.A2(n13769),
.A1(n11817),
.ZN(n11818));
NAND2_X1 U7763 (.A2(n11818),
.A1(n13782),
.ZN(n13846));
INV_X1 U7764 (.A(n13488),
.ZN(n12452));
NAND2_X1 U7765 (.A2(n12452),
.A1(n13782),
.ZN(n11819));
NAND2_X1 U7767 (.A2(n13785),
.A1(n13210),
.ZN(n11824));
AOI22_X1 U7768 (.B2(n11157),
.B1(REG2_REG_29__SCAN_IN),
.A1(FE_OFN8_n11821),
.A2(n11822),
.ZN(n11823));
OAI211_X1 U7769 (.C1(n13779),
.A(KgXiNKYImGwoITNkFdnqdBmiQCHYgIoS_ZN),
.C2(n11825),
.B(n11823),
.ZN(n11826));
NAND4_X1 U7770 (.A4(n11827),
.A3(n11828),
.A1(n11830),
.A2(n11829),
.ZN(U3354));
AOI22_X1 U7771 (.B2(n12169),
.B1(IR_REG_0__SCAN_IN),
.A1(FE_OFN0_n11847),
.A2(n12429),
.ZN(n11833));
NAND2_X1 U7772 (.A2(n11831),
.A1(FE_OFN0_n11847),
.ZN(n11837));
NAND2_X1 U7773 (.A2(REG1_REG_0__SCAN_IN),
.A1(n12169),
.ZN(n11836));
NAND2_X1 U7774 (.A2(n12429),
.A1(n12925),
.ZN(n11835));
NAND3_X1 U7775 (.A3(n11835),
.A1(n11837),
.A2(n11836),
.ZN(n12264));
NAND2_X1 U7776 (.A2(n12264),
.A1(n12265),
.ZN(n12263));
INV_X1 U7777 (.A(n12264),
.ZN(n11839));
NAND2_X1 U7778 (.A2(n11358),
.A1(FE_OFN0_n11847),
.ZN(n11844));
NAND2_X1 U7779 (.A2(n11842),
.A1(n12925),
.ZN(n11843));
NAND2_X1 U7780 (.A2(n11843),
.A1(n11844),
.ZN(n11845));
XNOR2_X1 U7781 (.B(FE_OFN5_n12926),
.A(n11845),
.ZN(n12309));
NOR2_X1 U7782 (.A2(n12309),
.A1(n12310),
.ZN(n11852));
AND2_X1 U7783 (.A2(n11842),
.A1(FE_OFN0_n11847),
.ZN(n11848));
AOI21_X1 U7784 (.A(n11848),
.B2(n11358),
.B1(n11846),
.ZN(n12311));
AND2_X1 U7785 (.A2(n13132),
.A1(FE_OFN0_n11847),
.ZN(n11849));
AOI21_X1 U7786 (.A(n11849),
.B2(FE_OFN20_n11698),
.B1(n11846),
.ZN(n11851));
OAI211_X1 U7787 (.C1(n11852),
.A(n11851),
.C2(n12311),
.B(n11853),
.ZN(n12384));
AOI22_X1 U7788 (.B2(n13132),
.B1(n12925),
.A1(FE_OFN0_n11847),
.A2(FE_OFN20_n11698),
.ZN(n11850));
XNOR2_X1 U7789 (.B(n11975),
.A(n11850),
.ZN(n12387));
AND2_X1 U7790 (.A2(n12490),
.A1(FE_OFN0_n11847),
.ZN(n11855));
AOI21_X1 U7791 (.A(n11855),
.B2(n13784),
.B1(n11846),
.ZN(n12412));
INV_X1 U7792 (.A(n12412),
.ZN(n11859));
NAND2_X1 U7793 (.A2(n13784),
.A1(FE_OFN0_n11847),
.ZN(n11857));
NAND2_X1 U7794 (.A2(n12490),
.A1(n12925),
.ZN(n11856));
NAND2_X1 U7795 (.A2(n11856),
.A1(n11857),
.ZN(n11858));
XNOR2_X1 U7796 (.B(FE_OFN5_n12926),
.A(n11858),
.ZN(n12411));
AOI22_X1 U7797 (.B2(n13138),
.B1(n12925),
.A1(FE_OFN0_n11847),
.A2(n13221),
.ZN(n11860));
XNOR2_X1 U7798 (.B(n11975),
.A(n11860),
.ZN(n11867));
INV_X2 U7799 (.A(n11846),
.ZN(n11977));
OAI22_X1 U7800 (.B2(n11884),
.B1(n13135),
.A1(n11977),
.A2(n13818),
.ZN(n11866));
OR2_X1 U7801 (.A2(n11866),
.A1(n11867),
.ZN(n12536));
AOI22_X1 U7802 (.B2(n12543),
.B1(n12925),
.A1(FE_OFN0_n11847),
.A2(n13220),
.ZN(n11861));
XNOR2_X1 U7803 (.B(n11975),
.A(n11861),
.ZN(n11869));
OAI22_X1 U7804 (.B2(n11884),
.B1(n11795),
.A1(n11977),
.A2(n12618),
.ZN(n11868));
NAND2_X1 U7805 (.A2(n12538),
.A1(n12536),
.ZN(n12610));
AOI22_X1 U7806 (.B2(n12654),
.B1(n12925),
.A1(FE_OFN0_n11847),
.A2(n13218),
.ZN(n11862));
XNOR2_X1 U7807 (.B(n11975),
.A(n11862),
.ZN(n11874));
OAI22_X1 U7808 (.B2(n11884),
.B1(n11863),
.A1(n11977),
.A2(n12675),
.ZN(n11873));
OR2_X1 U7809 (.A2(n11873),
.A1(n11874),
.ZN(n12648));
AOI22_X1 U7810 (.B2(n12620),
.B1(n12925),
.A1(FE_OFN0_n11847),
.A2(n13219),
.ZN(n11864));
XNOR2_X1 U7811 (.B(n11975),
.A(n11864),
.ZN(n11872));
OAI22_X1 U7812 (.B2(n11865),
.B1(n11884),
.A1(n11977),
.A2(n12652),
.ZN(n11871));
INV_X1 U7813 (.A(n12645),
.ZN(n12615));
NAND2_X1 U7814 (.A2(n12615),
.A1(n12648),
.ZN(n11878));
NOR2_X1 U7815 (.A2(n11878),
.A1(n12610),
.ZN(n11880));
NAND2_X1 U7816 (.A2(n11866),
.A1(n11867),
.ZN(n12466));
INV_X1 U7817 (.A(n12466),
.ZN(n12535));
NAND2_X1 U7818 (.A2(n11868),
.A1(n11869),
.ZN(n12537));
INV_X1 U7819 (.A(n12537),
.ZN(n11870));
AOI21_X1 U7820 (.A(n11870),
.B2(n12535),
.B1(n12538),
.ZN(n12611));
NAND2_X1 U7821 (.A2(n11871),
.A1(n11872),
.ZN(n12644));
INV_X1 U7822 (.A(n12644),
.ZN(n11876));
NAND2_X1 U7823 (.A2(n11873),
.A1(n11874),
.ZN(n12647));
INV_X1 U7824 (.A(n12647),
.ZN(n11875));
AOI21_X1 U7825 (.A(n11875),
.B2(n11876),
.B1(n12648),
.ZN(n11877));
OAI21_X1 U7826 (.A(n11877),
.B2(n11878),
.B1(n12611),
.ZN(n11879));
AOI22_X1 U7827 (.B2(n12677),
.B1(FE_OFN22_n12925),
.A1(FE_OFN0_n11847),
.A2(n13217),
.ZN(n11881));
XNOR2_X1 U7828 (.B(n11975),
.A(n11881),
.ZN(n11886));
OAI22_X1 U7829 (.B2(n12629),
.B1(n11884),
.A1(n11977),
.A2(n12828),
.ZN(n11885));
OR2_X1 U7830 (.A2(n11885),
.A1(n11886),
.ZN(n12749));
AOI22_X1 U7831 (.B2(n12757),
.B1(FE_OFN22_n12925),
.A1(FE_OFN0_n11847),
.A2(n13216),
.ZN(n11882));
XNOR2_X1 U7832 (.B(n11975),
.A(n11882),
.ZN(n11888));
OAI22_X1 U7833 (.B2(n11884),
.B1(n12827),
.A1(n11977),
.A2(n12794),
.ZN(n11887));
OR2_X1 U7834 (.A2(n11887),
.A1(n11888),
.ZN(n12752));
NAND2_X1 U7835 (.A2(n12752),
.A1(n12749),
.ZN(n12732));
AOI22_X1 U7836 (.B2(n12796),
.B1(FE_OFN22_n12925),
.A1(FE_OFN0_n11847),
.A2(n13215),
.ZN(n11883));
XNOR2_X1 U7837 (.B(n11975),
.A(n11883),
.ZN(n11891));
OAI22_X1 U7838 (.B2(n11884),
.B1(n12718),
.A1(n11977),
.A2(n13700),
.ZN(n11890));
NOR2_X1 U7839 (.A2(n11890),
.A1(n11891),
.ZN(n12736));
NAND2_X1 U7840 (.A2(n11885),
.A1(n11886),
.ZN(n12672));
INV_X1 U7841 (.A(n12672),
.ZN(n12748));
NAND2_X1 U7842 (.A2(n11887),
.A1(n11888),
.ZN(n12751));
INV_X1 U7843 (.A(n12751),
.ZN(n11889));
AOI21_X1 U7844 (.A(n11889),
.B2(n12748),
.B1(n12752),
.ZN(n12733));
NAND2_X1 U7845 (.A2(n11890),
.A1(n11891),
.ZN(n12737));
OAI21_X1 U7846 (.A(n12737),
.B2(n12736),
.B1(n12733),
.ZN(n11892));
INV_X1 U7847 (.A(n11892),
.ZN(n11893));
AOI22_X1 U7848 (.B2(n12822),
.B1(FE_OFN22_n12925),
.A1(FE_OFN0_n11847),
.A2(n13687),
.ZN(n11894));
XNOR2_X1 U7849 (.B(FE_OFN5_n12926),
.A(n11894),
.ZN(n12600));
AOI22_X1 U7850 (.B2(n12822),
.B1(FE_OFN0_n11847),
.A1(n11846),
.A2(n13687),
.ZN(n12601));
AOI22_X1 U7851 (.B2(n13572),
.B1(FE_OFN22_n12925),
.A1(FE_OFN0_n11847),
.A2(n13214),
.ZN(n11895));
XNOR2_X1 U7852 (.B(FE_OFN5_n12926),
.A(n11895),
.ZN(n12785));
AND2_X1 U7854 (.A2(n13572),
.A1(FE_OFN0_n11847),
.ZN(n11896));
AOI21_X1 U7855 (.A(n11896),
.B2(n13214),
.B1(n11846),
.ZN(n12784));
AND2_X1 U7856 (.A2(n13554),
.A1(FE_OFN0_n11847),
.ZN(n11902));
AOI21_X1 U7857 (.A(n11902),
.B2(n13689),
.B1(n11846),
.ZN(n11907));
NAND2_X1 U7858 (.A2(n13689),
.A1(FE_OFN0_n11847),
.ZN(n11904));
NAND2_X1 U7859 (.A2(n13554),
.A1(FE_OFN22_n12925),
.ZN(n11903));
NAND2_X1 U7860 (.A2(n11903),
.A1(n11904),
.ZN(n11905));
XNOR2_X1 U7861 (.B(n11975),
.A(n11905),
.ZN(n11906));
NOR2_X1 U7862 (.A2(n11906),
.A1(n11907),
.ZN(n12997));
INV_X1 U7863 (.A(n12997),
.ZN(n11908));
AND2_X1 U7864 (.A2(n11906),
.A1(n11907),
.ZN(n12996));
AOI22_X1 U7865 (.B2(FE_OFN22_n12925),
.B1(n13036),
.A1(n13655),
.A2(FE_OFN0_n11847),
.ZN(n11909));
XNOR2_X1 U7866 (.B(n11975),
.A(n11909),
.ZN(n11919));
OAI22_X1 U7867 (.B2(n11884),
.B1(n13670),
.A1(n11977),
.A2(n13526),
.ZN(n11918));
AOI22_X1 U7868 (.B2(n13534),
.B1(FE_OFN22_n12925),
.A1(n13666),
.A2(FE_OFN0_n11847),
.ZN(n11910));
XNOR2_X1 U7869 (.B(n11975),
.A(n11910),
.ZN(n11917));
OAI22_X1 U7870 (.B2(n11884),
.B1(n11911),
.A1(n11977),
.A2(n13545),
.ZN(n11916));
OR2_X1 U7871 (.A2(n11916),
.A1(n11917),
.ZN(n13029));
NAND2_X1 U7872 (.A2(n13029),
.A1(n11172),
.ZN(n12954));
AOI22_X1 U7873 (.B2(FE_OFN22_n12925),
.B1(FzxTCFmmmorPYWBoKVOYVzYHHyJMkxJR_ZN),
.A1(FE_OFN6_n13667),
.A2(FE_OFN0_n11847),
.ZN(n11912));
XNOR2_X1 U7874 (.B(n11975),
.A(n11912),
.ZN(n11922));
INV_X1 U7875 (.A(FE_OFN6_n13667),
.ZN(n11913));
OAI22_X1 U7876 (.B2(n11884),
.B1(n13658),
.A1(n11977),
.A2(n11913),
.ZN(n11921));
NOR2_X1 U7877 (.A2(n11921),
.A1(n11922),
.ZN(n12958));
NOR2_X1 U7878 (.A2(n12958),
.A1(n12954),
.ZN(n12971));
AOI22_X1 U7879 (.B2(n12976),
.B1(FE_OFN22_n12925),
.A1(n13656),
.A2(FE_OFN0_n11847),
.ZN(n11914));
XNOR2_X1 U7880 (.B(n11975),
.A(n11914),
.ZN(n11924));
OAI22_X1 U7881 (.B2(n13471),
.B1(n11884),
.A1(n11977),
.A2(n11915),
.ZN(n11923));
OR2_X1 U7882 (.A2(n11923),
.A1(n11924),
.ZN(n12973));
AND2_X1 U7883 (.A2(n12973),
.A1(n12971),
.ZN(n11928));
NAND2_X1 U7884 (.A2(n11916),
.A1(n11917),
.ZN(n12898));
INV_X1 U7885 (.A(n12898),
.ZN(n13028));
NAND2_X1 U7886 (.A2(n11918),
.A1(n11919),
.ZN(n13031));
INV_X1 U7887 (.A(n13031),
.ZN(n11920));
AOI21_X1 U7888 (.A(n11920),
.B2(n13028),
.B1(n11172),
.ZN(n12955));
NAND2_X1 U7889 (.A2(n11921),
.A1(n11922),
.ZN(n12959));
OAI21_X1 U7890 (.A(n12959),
.B2(n12958),
.B1(n12955),
.ZN(n12970));
NAND2_X1 U7891 (.A2(n11923),
.A1(n11924),
.ZN(n12972));
INV_X1 U7892 (.A(n12972),
.ZN(n11925));
AOI21_X1 U7893 (.A(n11925),
.B2(n12973),
.B1(n12970),
.ZN(n11926));
INV_X1 U7894 (.A(n11926),
.ZN(n11927));
AOI21_X1 U7895 (.A(n11927),
.B2(n11928),
.B1(n13030),
.ZN(n11930));
INV_X1 U7896 (.A(n11930),
.ZN(n13022));
AOI22_X1 U7897 (.B2(n13452),
.B1(FE_OFN22_n12925),
.A1(n13464),
.A2(FE_OFN0_n11847),
.ZN(n11929));
XNOR2_X1 U7898 (.B(FE_OFN5_n12926),
.A(n11929),
.ZN(n13020));
INV_X1 U7899 (.A(n13020),
.ZN(n11932));
AOI22_X1 U7900 (.B2(n13452),
.B1(FE_OFN0_n11847),
.A1(n11846),
.A2(n13464),
.ZN(n13019));
AOI21_X1 U7901 (.A(n13019),
.B2(n13020),
.B1(n11930),
.ZN(n11931));
AOI21_X1 U7902 (.A(n11931),
.B2(n11932),
.B1(n13022),
.ZN(n12942));
NAND2_X1 U7903 (.A2(FE_OFN0_n11847),
.A1(n13640),
.ZN(n11934));
NAND2_X1 U7904 (.A2(FE_OFN22_n12925),
.A1(n13438),
.ZN(n11933));
NAND2_X1 U7905 (.A2(n11933),
.A1(n11934),
.ZN(n11935));
XNOR2_X1 U7906 (.B(FE_OFN5_n12926),
.A(n11935),
.ZN(n12907));
NAND2_X1 U7910 (.A2(n12908),
.A1(n12907),
.ZN(n12940));
NAND2_X1 U7911 (.A2(FE_OFN0_n11847),
.A1(n13612),
.ZN(n11939));
NAND2_X1 U7912 (.A2(n13624),
.A1(FE_OFN22_n12925),
.ZN(n11938));
NAND2_X1 U7913 (.A2(n11938),
.A1(n11939),
.ZN(n11940));
XNOR2_X1 U7914 (.B(FE_OFN5_n12926),
.A(n11940),
.ZN(n12982));
NAND2_X1 U7916 (.A2(n11846),
.A1(n13612),
.ZN(n11942));
NAND2_X1 U7917 (.A2(n13624),
.A1(FE_OFN0_n11847),
.ZN(n11941));
NOR2_X1 U7920 (.A2(n12908),
.A1(n12907),
.ZN(n12941));
NAND2_X1 U7922 (.A2(FE_OFN0_n11847),
.A1(n13605),
.ZN(n11947));
NAND2_X1 U7923 (.A2(n13611),
.A1(FE_OFN22_n12925),
.ZN(n11946));
NAND2_X1 U7924 (.A2(n11946),
.A1(n11947),
.ZN(n11948));
XNOR2_X1 U7925 (.B(n11975),
.A(n11948),
.ZN(n11954));
AND2_X1 U7927 (.A2(n13611),
.A1(FE_OFN0_n11847),
.ZN(n11950));
AOI21_X1 U7928 (.A(n11950),
.B2(n11846),
.B1(n13605),
.ZN(n11953));
NAND2_X1 U7931 (.A2(n11953),
.A1(n11954),
.ZN(n12945));
INV_X1 U7932 (.A(n12945),
.ZN(n11955));
AOI22_X1 U7933 (.B2(n12889),
.B1(FE_OFN22_n12925),
.A1(n13343),
.A2(FE_OFN0_n11847),
.ZN(n11956));
XNOR2_X1 U7934 (.B(n11975),
.A(n11956),
.ZN(n11969));
OAI22_X1 U7935 (.B2(n12141),
.B1(n11884),
.A1(n13890),
.A2(n11977),
.ZN(n11968));
NOR2_X1 U7936 (.A2(n11968),
.A1(n11969),
.ZN(n12059));
AOI22_X1 U7937 (.B2(n13586),
.B1(FE_OFN22_n12925),
.A1(n13213),
.A2(FE_OFN0_n11847),
.ZN(n11957));
XNOR2_X1 U7938 (.B(n11975),
.A(n11957),
.ZN(n11967));
OAI22_X1 U7939 (.B2(n13337),
.B1(n11884),
.A1(n13355),
.A2(n11977),
.ZN(n11966));
NOR2_X1 U7940 (.A2(n11966),
.A1(n11967),
.ZN(n12103));
NOR2_X1 U7941 (.A2(n12103),
.A1(n12059),
.ZN(n11971));
AOI22_X1 U7942 (.B2(n13604),
.B1(FE_OFN22_n12925),
.A1(n13362),
.A2(FE_OFN0_n11847),
.ZN(n11958));
XNOR2_X1 U7943 (.B(n11975),
.A(n11958),
.ZN(n11963));
OAI22_X1 U7944 (.B2(n13384),
.B1(n11884),
.A1(n13614),
.A2(n11977),
.ZN(n11962));
NOR2_X1 U7945 (.A2(n11962),
.A1(n11963),
.ZN(n12072));
AOI22_X1 U7946 (.B2(n13360),
.B1(FE_OFN22_n12925),
.A1(n13587),
.A2(FE_OFN0_n11847),
.ZN(n11960));
XNOR2_X1 U7947 (.B(n11975),
.A(n11960),
.ZN(n11965));
OAI22_X1 U7948 (.B2(n13595),
.B1(n11884),
.A1(n13341),
.A2(n11977),
.ZN(n11964));
NOR2_X1 U7949 (.A2(n11964),
.A1(n11965),
.ZN(n12074));
NOR2_X1 U7950 (.A2(n12074),
.A1(n12072),
.ZN(n12102));
NAND2_X1 U7951 (.A2(n12102),
.A1(n11971),
.ZN(n12086));
AOI22_X1 U7952 (.B2(n12877),
.B1(FE_OFN22_n12925),
.A1(n13212),
.A2(FE_OFN0_n11847),
.ZN(n11961));
XNOR2_X1 U7953 (.B(n11975),
.A(n11961),
.ZN(n11973));
INV_X1 U7954 (.A(n13212),
.ZN(n12132));
OAI22_X1 U7955 (.B2(n12032),
.B1(n11884),
.A1(n12132),
.A2(n11977),
.ZN(n11972));
NOR2_X1 U7956 (.A2(n11972),
.A1(n11973),
.ZN(n12090));
NOR2_X1 U7957 (.A2(n12090),
.A1(n12086),
.ZN(n12917));
NAND2_X1 U7958 (.A2(n11962),
.A1(n11963),
.ZN(n13007));
NAND2_X1 U7959 (.A2(n11964),
.A1(n11965),
.ZN(n12075));
OAI21_X1 U7960 (.A(n12075),
.B2(n13007),
.B1(n12074),
.ZN(n12101));
NAND2_X1 U7961 (.A2(n11966),
.A1(n11967),
.ZN(n12104));
NAND2_X1 U7962 (.A2(n11968),
.A1(n11969),
.ZN(n12060));
OAI21_X1 U7963 (.A(n12060),
.B2(n12104),
.B1(n12059),
.ZN(n11970));
AOI21_X1 U7964 (.A(n11970),
.B2(n12101),
.B1(n11971),
.ZN(n12087));
NAND2_X1 U7965 (.A2(n11972),
.A1(n11973),
.ZN(n12091));
OAI21_X1 U7966 (.A(n12091),
.B2(n12090),
.B1(n12087),
.ZN(n12920));
AOI21_X1 U7967 (.A(n12920),
.B2(n12917),
.B1(n13010),
.ZN(n11980));
AOI22_X1 U7968 (.B2(n11974),
.B1(FE_OFN22_n12925),
.A1(n13211),
.A2(FE_OFN0_n11847),
.ZN(n11976));
XNOR2_X1 U7969 (.B(n11975),
.A(n11976),
.ZN(n11979));
OAI22_X1 U7970 (.B2(n13324),
.B1(n11884),
.A1(n12935),
.A2(n11977),
.ZN(n11978));
NAND2_X1 U7971 (.A2(n11978),
.A1(n11979),
.ZN(n12918));
XNOR2_X1 U7972 (.B(n11309),
.A(n11980),
.ZN(n11988));
NAND2_X1 U7973 (.A2(n11982),
.A1(n11983),
.ZN(n11987));
NAND3_X1 U7974 (.A3(n11984),
.A1(n11986),
.A2(n11985),
.ZN(n11989));
NAND2_X1 U7975 (.A2(n11997),
.A1(n11987),
.ZN(n13005));
NAND2_X1 U7976 (.A2(n13043),
.A1(n11988),
.ZN(n12001));
NAND2_X1 U7977 (.A2(n11989),
.A1(n11990),
.ZN(n11991));
NAND2_X1 U7978 (.A2(n13203),
.A1(n11991),
.ZN(n12315));
OAI21_X1 U7979 (.A(STATE_REG_SCAN_IN),
.B2(n12169),
.B1(n12315),
.ZN(n11992));
OR2_X1 U7980 (.A2(U3149),
.A1(n12170),
.ZN(n13815));
NAND2_X1 U7981 (.A2(n13623),
.A1(n11997),
.ZN(n11993));
OAI22_X1 U7982 (.B2(n11994),
.B1(STATE_REG_SCAN_IN),
.A1(n12991),
.A2(n13324),
.ZN(n11996));
NAND3_X2 U7983 (.A3(n13203),
.A1(n11997),
.A2(n13688),
.ZN(n12990));
NOR2_X1 U7984 (.A2(n12990),
.A1(n12132),
.ZN(n11995));
AOI211_X1 U7985 (.C1(n13328),
.A(n11996),
.C2(n13016),
.B(n11995),
.ZN(n11999));
NAND2_X1 U7986 (.A2(n12000),
.A1(n12001),
.ZN(U3211));
NAND2_X1 U7987 (.A2(n13672),
.A1(n12120),
.ZN(n12010));
INV_X1 U7988 (.A(n13209),
.ZN(n12008));
AOI22_X1 U7989 (.B2(n13623),
.B1(n12932),
.A1(n13211),
.A2(n13688),
.ZN(n12007));
OAI21_X1 U7990 (.A(n12007),
.B2(n13627),
.B1(n12008),
.ZN(n12009));
INV_X1 U7992 (.A(n12011),
.ZN(n12051));
OR2_X2 U7996 (.A2(n12124),
.A1(n12127),
.ZN(n12129));
XNOR2_X1 U7997 (.B(n12877),
.A(n13212),
.ZN(n13117));
NAND2_X1 U7998 (.A2(n12019),
.A1(n12130),
.ZN(n12021));
NAND2_X1 U7999 (.A2(n12020),
.A1(n12021),
.ZN(n12022));
XNOR2_X1 U8000 (.B(n13117),
.A(n12022),
.ZN(n12885));
NOR2_X1 U8001 (.A2(n12032),
.A1(n13698),
.ZN(n12023));
AOI21_X1 U8002 (.A(n12023),
.B2(n13688),
.B1(n13343),
.ZN(n12024));
OAI21_X1 U8003 (.A(n12024),
.B2(n13627),
.B1(n12935),
.ZN(n12025));
AOI21_X1 U8004 (.A(n12025),
.B2(n13672),
.B1(n12885),
.ZN(n12026));
MUX2_X1 U8005 (.S(n13839),
.A(n12035),
.B(REG1_REG_26__SCAN_IN),
.Z(n12029));
INV_X1 U8006 (.A(n12029),
.ZN(n12034));
OAI21_X1 U8007 (.A(n12031),
.B2(n12032),
.B1(n12030),
.ZN(n12883));
NAND2_X1 U8008 (.A2(n13374),
.A1(n13841),
.ZN(n13835));
NAND2_X1 U8009 (.A2(n12033),
.A1(n12034),
.ZN(U3544));
MUX2_X1 U8010 (.S(FE_OFN3_n13832),
.A(REG0_REG_26__SCAN_IN),
.B(n12035),
.Z(n12036));
INV_X1 U8011 (.A(n12036),
.ZN(n12038));
NAND2_X1 U8012 (.A2(n12037),
.A1(n12038),
.ZN(U3512));
XNOR2_X1 U8013 (.B(n13113),
.A(n12041),
.ZN(n13322));
XNOR2_X1 U8014 (.B(n13113),
.A(n12042),
.ZN(n12046));
OAI21_X1 U8015 (.A(n13331),
.B2(n13698),
.B1(n13324),
.ZN(n12047));
NAND2_X1 U8016 (.A2(FE_OFN3_n13832),
.A1(n12149),
.ZN(n12050));
INV_X1 U8017 (.A(REG0_REG_27__SCAN_IN),
.ZN(n12048));
NAND2_X1 U8018 (.A2(n12048),
.A1(n13860),
.ZN(n12049));
NAND2_X1 U8019 (.A2(n12049),
.A1(n12050),
.ZN(n12054));
INV_X1 U8020 (.A(n12031),
.ZN(n12052));
OR2_X1 U8021 (.A2(FE_OFN21_n13759),
.A1(n13325),
.ZN(n12053));
NAND2_X1 U8022 (.A2(n12053),
.A1(n12054),
.ZN(U3513));
INV_X1 U8023 (.A(n12102),
.ZN(n12055));
NOR2_X1 U8024 (.A2(n12103),
.A1(n12055),
.ZN(n12058));
INV_X1 U8025 (.A(n12101),
.ZN(n12056));
OAI21_X1 U8026 (.A(n12104),
.B2(n12103),
.B1(n12056),
.ZN(n12057));
AOI21_X1 U8027 (.A(n12057),
.B2(n12058),
.B1(n13010),
.ZN(n12062));
XNOR2_X1 U8029 (.B(n11311),
.A(n12062),
.ZN(n12063));
NAND2_X1 U8030 (.A2(n13043),
.A1(n12063),
.ZN(n12071));
INV_X1 U8031 (.A(n12064),
.ZN(n12891));
AOI22_X1 U8032 (.B2(U3149),
.B1(REG3_REG_25__SCAN_IN),
.A1(n13037),
.A2(n12889),
.ZN(n12065));
OAI21_X1 U8033 (.A(n12065),
.B2(n13041),
.B1(n12891),
.ZN(n12066));
AOI21_X1 U8034 (.A(n12066),
.B2(n13213),
.B1(n13038),
.ZN(n12067));
NAND2_X1 U8036 (.A2(n12070),
.A1(n12071),
.ZN(U3222));
INV_X1 U8037 (.A(n12072),
.ZN(n13008));
INV_X1 U8038 (.A(n13007),
.ZN(n12073));
AOI21_X1 U8039 (.A(n12073),
.B2(n13008),
.B1(n13010),
.ZN(n12077));
XNOR2_X1 U8041 (.B(n11303),
.A(n12077),
.ZN(n12078));
NAND2_X1 U8042 (.A2(n13043),
.A1(n12078),
.ZN(n12085));
INV_X1 U8043 (.A(n12079),
.ZN(n13361));
AOI22_X1 U8044 (.B2(U3149),
.B1(REG3_REG_23__SCAN_IN),
.A1(n13362),
.A2(n13038),
.ZN(n12080));
OAI21_X1 U8045 (.A(n12080),
.B2(n13595),
.B1(n12991),
.ZN(n12081));
NAND2_X1 U8048 (.A2(n12084),
.A1(n12085),
.ZN(U3213));
INV_X1 U8049 (.A(n12086),
.ZN(n12089));
INV_X1 U8050 (.A(n12087),
.ZN(n12088));
AOI21_X1 U8051 (.A(n12088),
.B2(n12089),
.B1(n13010),
.ZN(n12093));
XNOR2_X1 U8053 (.B(n11310),
.A(n12093),
.ZN(n12094));
NAND2_X1 U8054 (.A2(n13043),
.A1(n12094),
.ZN(n12100));
AOI22_X1 U8055 (.B2(U3149),
.B1(REG3_REG_26__SCAN_IN),
.A1(n13037),
.A2(n12877),
.ZN(n12095));
OAI21_X1 U8056 (.A(n12095),
.B2(n13041),
.B1(n12880),
.ZN(n12096));
AOI21_X1 U8057 (.A(n12096),
.B2(n13343),
.B1(n13038),
.ZN(n12097));
NAND2_X1 U8058 (.A2(n12099),
.A1(n12100),
.ZN(U3237));
XNOR2_X1 U8060 (.B(n11312),
.A(n12106),
.ZN(n12107));
NAND2_X1 U8061 (.A2(n13043),
.A1(n12107),
.ZN(n12113));
AOI22_X1 U8062 (.B2(U3149),
.B1(REG3_REG_24__SCAN_IN),
.A1(n13037),
.A2(n13586),
.ZN(n12108));
OAI21_X1 U8063 (.A(n12108),
.B2(n12990),
.B1(n13341),
.ZN(n12109));
AOI21_X1 U8064 (.A(n12109),
.B2(n13016),
.B1(n13338),
.ZN(n12110));
OAI21_X1 U8065 (.A(n12110),
.B2(n13014),
.B1(n13890),
.ZN(n12111));
INV_X1 U8066 (.A(n12111),
.ZN(n12112));
NAND2_X1 U8067 (.A2(n12112),
.A1(n12113),
.ZN(U3226));
NOR2_X1 U8068 (.A2(n13627),
.A1(n11157),
.ZN(n13571));
NAND2_X1 U8069 (.A2(n13785),
.A1(n13211),
.ZN(n12115));
AOI22_X1 U8070 (.B2(n11157),
.B1(REG2_REG_28__SCAN_IN),
.A1(FE_OFN8_n11821),
.A2(n12932),
.ZN(n12114));
OAI211_X1 U8071 (.C1(n13779),
.A(n12115),
.C2(n12934),
.B(n12114),
.ZN(n12397));
AOI21_X1 U8072 (.A(n12116),
.B2(n13209),
.B1(FE_OFN10_n13571),
.ZN(n12117));
NOR2_X1 U8074 (.A2(n13568),
.A1(n11157),
.ZN(n13503));
NOR2_X1 U8075 (.A2(n13584),
.A1(n12118),
.ZN(n12119));
NAND2_X1 U8079 (.A2(n12125),
.A1(n12126),
.ZN(n13071));
INV_X1 U8080 (.A(n12135),
.ZN(n12897));
OAI22_X1 U8081 (.B2(n13698),
.B1(n12141),
.A1(n13355),
.A2(n13819),
.ZN(n13907));
NAND2_X1 U8082 (.A2(n13072),
.A1(n12130),
.ZN(n12131));
XNOR2_X1 U8083 (.B(n13071),
.A(n12131),
.ZN(n12133));
OAI21_X1 U8086 (.A(n12140),
.B2(n12141),
.B1(n12139),
.ZN(n12892));
NAND2_X1 U8087 (.A2(REG0_REG_25__SCAN_IN),
.A1(n13860),
.ZN(n12142));
NAND2_X1 U8090 (.A2(n13841),
.A1(n12160),
.ZN(n12165));
NAND2_X1 U8091 (.A2(REG1_REG_29__SCAN_IN),
.A1(n13839),
.ZN(n12161));
INV_X1 U8092 (.A(n12163),
.ZN(n12164));
NAND2_X1 U8093 (.A2(n12164),
.A1(n12165),
.ZN(U3547));
NOR2_X1 U8094 (.A2(U3149),
.A1(n12166),
.ZN(n12167));
NAND2_X1 U8097 (.A2(n12169),
.A1(n12170),
.ZN(n12171));
NAND2_X1 U8098 (.A2(STATE_REG_SCAN_IN),
.A1(n12171),
.ZN(n12189));
NOR2_X1 U8100 (.A2(n11687),
.A1(n11686),
.ZN(n12174));
NAND3_X1 U8101 (.A3(REG2_REG_0__SCAN_IN),
.A1(IR_REG_0__SCAN_IN),
.A2(REG2_REG_1__SCAN_IN),
.ZN(n12297));
AOI21_X1 U8102 (.A(REG2_REG_1__SCAN_IN),
.B2(REG2_REG_0__SCAN_IN),
.B1(IR_REG_0__SCAN_IN),
.ZN(n12299));
NAND2_X1 U8103 (.A2(REG2_REG_2__SCAN_IN),
.A1(n12175),
.ZN(n13228));
NAND2_X1 U8104 (.A2(n13777),
.A1(n13228),
.ZN(n12178));
NAND3_X1 U8108 (.A3(n12240),
.A1(n13798),
.A2(n12498),
.ZN(n12184));
INV_X1 U8109 (.A(n12227),
.ZN(n12182));
NAND3_X1 U8111 (.A3(REG1_REG_0__SCAN_IN),
.A1(IR_REG_0__SCAN_IN),
.A2(REG1_REG_1__SCAN_IN),
.ZN(n12294));
AOI21_X1 U8112 (.A(REG1_REG_1__SCAN_IN),
.B2(REG1_REG_0__SCAN_IN),
.B1(IR_REG_0__SCAN_IN),
.ZN(n12296));
NAND2_X1 U8113 (.A2(REG1_REG_2__SCAN_IN),
.A1(n12179),
.ZN(n13226));
INV_X1 U8115 (.A(REG1_REG_2__SCAN_IN),
.ZN(n12454));
NAND2_X1 U8116 (.A2(n12441),
.A1(n12181),
.ZN(n12250));
NAND2_X1 U8117 (.A2(n12250),
.A1(n12249),
.ZN(n12185));
NAND2_X1 U8118 (.A2(n12185),
.A1(n13804),
.ZN(n12183));
NAND3_X1 U8119 (.A3(n13801),
.A1(n12184),
.A2(n12183),
.ZN(n12188));
OAI22_X1 U8121 (.B2(n12185),
.B1(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.A1(n13795),
.A2(n12186),
.ZN(n12187));
MUX2_X1 U8123 (.S(n12248),
.A(n12188),
.B(n12187),
.Z(n12194));
NAND2_X1 U8124 (.A2(REG2_REG_3__SCAN_IN),
.A1(n13776),
.ZN(n12243));
NOR3_X1 U8125 (.A3(n12243),
.A1(n13795),
.A2(n12240),
.ZN(n12193));
INV_X1 U8126 (.A(REG3_REG_3__SCAN_IN),
.ZN(n12413));
NOR2_X1 U8127 (.A2(n12413),
.A1(STATE_REG_SCAN_IN),
.ZN(n12192));
AOI21_X1 U8128 (.A(n12189),
.B2(n11569),
.B1(n12190),
.ZN(n13320));
AND2_X1 U8129 (.A2(ADDR_REG_3__SCAN_IN),
.A1(FE_OFN1_n13320),
.ZN(n12191));
OR4_X1 U8130 (.A4(n12191),
.A3(n12192),
.A1(n12194),
.A2(n12193),
.ZN(U3243));
MUX2_X1 U8131 (.S(U3149),
.A(n12379),
.B(n11432),
.Z(n12195));
INV_X1 U8132 (.A(n12195),
.ZN(U3345));
INV_X1 U8133 (.A(n12196),
.ZN(n12200));
NOR2_X1 U8134 (.A2(n12198),
.A1(U3149),
.ZN(n12839));
NAND2_X1 U8135 (.A2(n12839),
.A1(n12197),
.ZN(n12207));
AOI22_X1 U8137 (.B2(U3149),
.B1(DATAI_24_),
.A1(n12214),
.A2(IR_REG_24__SCAN_IN),
.ZN(n12199));
OAI21_X1 U8138 (.A(n12199),
.B2(n12207),
.B1(n12200),
.ZN(U3328));
NAND3_X1 U8140 (.A3(n12201),
.A1(n11495),
.A2(n12839),
.ZN(n12203));
NAND2_X1 U8141 (.A2(U3149),
.A1(DATAI_8_),
.ZN(n12202));
OAI211_X1 U8142 (.C1(n11447),
.A(n12203),
.C2(n12204),
.B(n12202),
.ZN(U3344));
INV_X1 U8143 (.A(DATAI_4_),
.ZN(n12205));
INV_X1 U8144 (.A(n12252),
.ZN(n12277));
MUX2_X1 U8145 (.S(STATE_REG_SCAN_IN),
.A(n12205),
.B(n12277),
.Z(n12206));
INV_X1 U8146 (.A(n12206),
.ZN(U3348));
INV_X1 U8147 (.A(DATAI_25_),
.ZN(n12210));
NAND2_X1 U8148 (.A2(STATE_REG_SCAN_IN),
.A1(n11758),
.ZN(n12208));
MUX2_X1 U8149 (.S(n11329),
.A(n12208),
.B(n12207),
.Z(n12209));
OAI21_X1 U8150 (.A(n12209),
.B2(n12210),
.B1(STATE_REG_SCAN_IN),
.ZN(U3327));
MUX2_X1 U8151 (.S(STATE_REG_SCAN_IN),
.A(n11497),
.B(n13269),
.Z(n12211));
INV_X1 U8152 (.A(n12211),
.ZN(U3339));
NAND3_X1 U8153 (.A3(n12212),
.A1(n12213),
.A2(n12839),
.ZN(n12216));
AOI22_X1 U8154 (.B2(U3149),
.B1(DATAI_18_),
.A1(n12214),
.A2(IR_REG_18__SCAN_IN),
.ZN(n12215));
NAND2_X1 U8155 (.A2(n12215),
.A1(n12216),
.ZN(U3334));
MUX2_X1 U8156 (.S(U3149),
.A(n13288),
.B(n11515),
.Z(n12217));
INV_X1 U8157 (.A(n12217),
.ZN(U3336));
INV_X1 U8158 (.A(DATAI_12_),
.ZN(n12218));
INV_X1 U8159 (.A(n12575),
.ZN(n13257));
MUX2_X1 U8160 (.S(STATE_REG_SCAN_IN),
.A(n12218),
.B(n13257),
.Z(n12219));
INV_X1 U8161 (.A(n12219),
.ZN(U3340));
INV_X1 U8162 (.A(DATAI_15_),
.ZN(n12220));
INV_X1 U8163 (.A(n12766),
.ZN(n12773));
MUX2_X1 U8164 (.S(STATE_REG_SCAN_IN),
.A(n12220),
.B(n12773),
.Z(n12221));
INV_X1 U8165 (.A(n12221),
.ZN(U3337));
INV_X1 U8166 (.A(D_REG_0__SCAN_IN),
.ZN(n12225));
INV_X1 U8167 (.A(n12223),
.ZN(n12224));
AOI22_X1 U8168 (.B2(n13204),
.B1(n12224),
.A1(n13814),
.A2(n12225),
.ZN(U3458));
NAND2_X1 U8169 (.A2(DATAO_REG_30__SCAN_IN),
.A1(n13223),
.ZN(n12226));
OAI21_X1 U8170 (.A(n12226),
.B2(n13223),
.B1(n13197),
.ZN(U3580));
INV_X1 U8171 (.A(REG3_REG_0__SCAN_IN),
.ZN(n12550));
AOI21_X1 U8172 (.A(IR_REG_0__SCAN_IN),
.B2(n11360),
.B1(n11687),
.ZN(n12229));
OAI21_X1 U8173 (.A(n13764),
.B2(REG2_REG_0__SCAN_IN),
.B1(n11687),
.ZN(n12228));
NAND2_X1 U8174 (.A2(n11236),
.A1(n12228),
.ZN(n12267));
OAI211_X1 U8175 (.C1(n12229),
.A(n12227),
.C2(n12228),
.B(n12267),
.ZN(n12230));
OAI21_X1 U8176 (.A(n12230),
.B2(n12550),
.B1(STATE_REG_SCAN_IN),
.ZN(n12232));
NOR3_X1 U8177 (.A3(n11236),
.A1(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.A2(REG1_REG_0__SCAN_IN),
.ZN(n12231));
AOI211_X1 U8178 (.C1(FE_OFN1_n13320),
.A(n12232),
.C2(ADDR_REG_0__SCAN_IN),
.B(n12231),
.ZN(n12233));
INV_X1 U8179 (.A(n12233),
.ZN(U3240));
NAND2_X1 U8180 (.A2(n11831),
.A1(n12863),
.ZN(n13124));
AOI22_X1 U8183 (.B2(n12429),
.B1(n12234),
.A1(n13690),
.A2(n11358),
.ZN(n12235));
OAI21_X1 U8184 (.A(n12235),
.B2(n13078),
.B1(n13619),
.ZN(n12236));
AOI21_X1 U8185 (.A(n12236),
.B2(n12237),
.B1(n13672),
.ZN(n13817));
NAND2_X1 U8186 (.A2(REG1_REG_0__SCAN_IN),
.A1(n13839),
.ZN(n12238));
OAI21_X1 U8187 (.A(n12238),
.B2(n13839),
.B1(n13817),
.ZN(U3518));
NOR2_X1 U8188 (.A2(U4043),
.A1(FE_OFN1_n13320),
.ZN(U3148));
NAND2_X1 U8189 (.A2(REG3_REG_5__SCAN_IN),
.A1(U3149),
.ZN(n12541));
INV_X1 U8190 (.A(n12541),
.ZN(n12261));
NAND2_X1 U8191 (.A2(n12243),
.A1(n12240),
.ZN(n12239));
NAND2_X1 U8192 (.A2(n12498),
.A1(n12248),
.ZN(n12241));
NAND3_X1 U8193 (.A3(REG2_REG_4__SCAN_IN),
.A1(n12239),
.A2(n12241),
.ZN(n12271));
NAND2_X1 U8194 (.A2(n12277),
.A1(n12271),
.ZN(n12246));
INV_X1 U8195 (.A(n12240),
.ZN(n12242));
NAND2_X1 U8199 (.A2(n12272),
.A1(n12246),
.ZN(n12247));
OR2_X1 U8200 (.A2(n11395),
.A1(n12247),
.ZN(n12286));
NAND2_X1 U8201 (.A2(n13580),
.A1(n12247),
.ZN(n12285));
NAND2_X1 U8202 (.A2(n12285),
.A1(n12286),
.ZN(n12255));
NAND2_X1 U8203 (.A2(n12250),
.A1(n12251),
.ZN(n12253));
INV_X1 U8204 (.A(REG1_REG_4__SCAN_IN),
.ZN(n12463));
XNOR2_X1 U8205 (.B(REG1_REG_5__SCAN_IN),
.A(n12283),
.ZN(n12254));
OAI22_X1 U8206 (.B2(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.B1(n12254),
.A1(n13795),
.A2(n12255),
.ZN(n12259));
INV_X1 U8207 (.A(n12254),
.ZN(n12257));
NAND2_X1 U8208 (.A2(n12255),
.A1(n13798),
.ZN(n12256));
OAI211_X1 U8209 (.C1(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.A(n12256),
.C2(n12257),
.B(n13801),
.ZN(n12258));
MUX2_X1 U8210 (.S(n13775),
.A(n12259),
.B(n12258),
.Z(n12260));
AOI211_X1 U8211 (.C1(FE_OFN1_n13320),
.A(n12261),
.C2(ADDR_REG_5__SCAN_IN),
.B(n12260),
.ZN(n12262));
INV_X1 U8212 (.A(n12262),
.ZN(U3245));
NAND2_X1 U8213 (.A2(REG2_REG_0__SCAN_IN),
.A1(IR_REG_0__SCAN_IN),
.ZN(n12266));
OAI21_X1 U8214 (.A(n12263),
.B2(n12264),
.B1(n12265),
.ZN(n12859));
MUX2_X1 U8215 (.S(n11687),
.A(n12266),
.B(n12859),
.Z(n12268));
OAI211_X1 U8216 (.C1(n12268),
.A(U4043),
.C2(n11686),
.B(n12267),
.ZN(n13238));
AND2_X1 U8217 (.A2(REG3_REG_4__SCAN_IN),
.A1(U3149),
.ZN(n12468));
NAND2_X1 U8218 (.A2(n12269),
.A1(n12270),
.ZN(n12275));
INV_X1 U8219 (.A(n12275),
.ZN(n12274));
NAND2_X1 U8220 (.A2(n12271),
.A1(n12272),
.ZN(n12276));
NAND2_X1 U8221 (.A2(n12276),
.A1(n13798),
.ZN(n12273));
OAI211_X1 U8222 (.C1(n12274),
.A(n12273),
.C2(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.B(n13801),
.ZN(n12279));
OAI22_X1 U8223 (.B2(n12275),
.B1(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.A1(n13795),
.A2(n12276),
.ZN(n12278));
MUX2_X1 U8224 (.S(n12277),
.A(n12279),
.B(n12278),
.Z(n12280));
AOI211_X1 U8225 (.C1(FE_OFN1_n13320),
.A(n12468),
.C2(ADDR_REG_4__SCAN_IN),
.B(n12280),
.ZN(n12281));
NAND2_X1 U8226 (.A2(n12281),
.A1(n13238),
.ZN(U3244));
AND2_X1 U8227 (.A2(REG1_REG_5__SCAN_IN),
.A1(n13775),
.ZN(n12282));
INV_X1 U8229 (.A(n12328),
.ZN(n13774));
XNOR2_X1 U8230 (.B(n13774),
.A(n12284),
.ZN(n12293));
NAND2_X1 U8231 (.A2(REG3_REG_6__SCAN_IN),
.A1(U3149),
.ZN(n12617));
INV_X1 U8232 (.A(n12617),
.ZN(n12291));
NAND2_X1 U8233 (.A2(n13775),
.A1(n12285),
.ZN(n12287));
NAND2_X1 U8234 (.A2(n12286),
.A1(n12287),
.ZN(n12330));
XNOR2_X1 U8235 (.B(REG2_REG_6__SCAN_IN),
.A(n12328),
.ZN(n12288));
XNOR2_X1 U8236 (.B(n12288),
.A(n12330),
.ZN(n12289));
OAI22_X1 U8237 (.B2(n13801),
.B1(n12328),
.A1(n13795),
.A2(n12289),
.ZN(n12290));
AOI211_X1 U8238 (.C1(FE_OFN1_n13320),
.A(n12291),
.C2(ADDR_REG_6__SCAN_IN),
.B(n12290),
.ZN(n12292));
OAI21_X1 U8239 (.A(n12292),
.B2(n12293),
.B1(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.ZN(U3246));
INV_X1 U8240 (.A(n12294),
.ZN(n12295));
NOR2_X1 U8241 (.A2(n12295),
.A1(n12296),
.ZN(n12304));
INV_X1 U8242 (.A(n12297),
.ZN(n12298));
NOR2_X1 U8243 (.A2(n12298),
.A1(n12299),
.ZN(n12303));
INV_X1 U8244 (.A(n12303),
.ZN(n12300));
NAND2_X1 U8245 (.A2(n12300),
.A1(n13798),
.ZN(n12301));
OAI211_X1 U8246 (.C1(n12304),
.A(n12301),
.C2(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.B(n13801),
.ZN(n12302));
INV_X1 U8247 (.A(n12302),
.ZN(n12306));
AOI22_X1 U8248 (.B2(n12303),
.B1(n13798),
.A1(n13804),
.A2(n12304),
.ZN(n12305));
AOI22_X1 U8249 (.B2(U3149),
.B1(REG3_REG_1__SCAN_IN),
.A1(FE_OFN1_n13320),
.A2(ADDR_REG_1__SCAN_IN),
.ZN(n12307));
NAND2_X1 U8250 (.A2(n12307),
.A1(n12308),
.ZN(U3241));
XOR2_X1 U8251 (.B(n12309),
.A(n12310),
.Z(n12313));
INV_X1 U8252 (.A(n12313),
.ZN(n12312));
MUX2_X1 U8253 (.S(n12311),
.A(n12313),
.B(n12312),
.Z(n12318));
AOI22_X1 U8254 (.B2(FE_OFN20_n11698),
.B1(n13035),
.A1(n13038),
.A2(n11831),
.ZN(n12317));
OR2_X1 U8255 (.A2(n12314),
.A1(n12315),
.ZN(n12860));
AOI22_X1 U8256 (.B2(n11842),
.B1(n13037),
.A1(n12860),
.A2(REG3_REG_1__SCAN_IN),
.ZN(n12316));
OAI211_X1 U8257 (.C1(n12318),
.A(n12317),
.C2(n13005),
.B(n12316),
.ZN(U3219));
NAND2_X1 U8258 (.A2(REG3_REG_8__SCAN_IN),
.A1(U3149),
.ZN(n12674));
INV_X1 U8259 (.A(n12674),
.ZN(n12346));
NAND2_X1 U8260 (.A2(n11409),
.A1(n12320),
.ZN(n12319));
NOR2_X1 U8263 (.A2(n12642),
.A1(n12379),
.ZN(n12325));
NAND2_X1 U8264 (.A2(n12642),
.A1(n12379),
.ZN(n12324));
AND2_X1 U8265 (.A2(REG1_REG_8__SCAN_IN),
.A1(n12324),
.ZN(n12323));
NAND3_X1 U8269 (.A3(n12349),
.A1(n13804),
.A2(n12348),
.ZN(n12339));
INV_X1 U8270 (.A(REG2_REG_6__SCAN_IN),
.ZN(n12508));
NAND2_X1 U8271 (.A2(n12508),
.A1(n12328),
.ZN(n12329));
NAND2_X1 U8275 (.A2(n12375),
.A1(n12379),
.ZN(n12333));
INV_X1 U8277 (.A(n12379),
.ZN(n12334));
XNOR2_X1 U8280 (.B(REG2_REG_8__SCAN_IN),
.A(n12356),
.ZN(n12340));
INV_X1 U8281 (.A(n12340),
.ZN(n12337));
NAND2_X1 U8282 (.A2(n12337),
.A1(n13798),
.ZN(n12338));
NAND2_X1 U8283 (.A2(n12338),
.A1(n12339),
.ZN(n12344));
AND2_X1 U8284 (.A2(n12349),
.A1(n12348),
.ZN(n12342));
NAND2_X1 U8285 (.A2(n12340),
.A1(n13798),
.ZN(n12341));
OAI211_X1 U8286 (.C1(n12342),
.A(n12341),
.C2(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.B(n13801),
.ZN(n12343));
MUX2_X1 U8287 (.S(n12357),
.A(n12344),
.B(n12343),
.Z(n12345));
AOI211_X1 U8288 (.C1(FE_OFN1_n13320),
.A(n12346),
.C2(ADDR_REG_8__SCAN_IN),
.B(n12345),
.ZN(n12347));
INV_X1 U8289 (.A(n12347),
.ZN(U3248));
NAND2_X1 U8290 (.A2(REG3_REG_9__SCAN_IN),
.A1(U3149),
.ZN(n12755));
INV_X1 U8291 (.A(n12755),
.ZN(n12370));
NAND2_X1 U8293 (.A2(WxUoeaFQeyYVaGStCqAbTWICyXpTFvtD_Z),
.A1(n12348),
.ZN(n12350));
NAND2_X1 U8294 (.A2(n12349),
.A1(n12350),
.ZN(n12351));
INV_X1 U8295 (.A(REG1_REG_9__SCAN_IN),
.ZN(n12835));
NAND2_X1 U8296 (.A2(n12835),
.A1(n12351),
.ZN(n12392));
INV_X1 U8297 (.A(n12351),
.ZN(n12352));
NAND3_X1 U8298 (.A3(n12393),
.A1(n13804),
.A2(n12392),
.ZN(n12362));
INV_X1 U8299 (.A(REG2_REG_8__SCAN_IN),
.ZN(n12353));
NAND2_X1 U8300 (.A2(n12353),
.A1(WxUoeaFQeyYVaGStCqAbTWICyXpTFvtD_Z),
.ZN(n12355));
NAND2_X1 U8301 (.A2(n12355),
.A1(n12356),
.ZN(n12359));
NAND2_X1 U8302 (.A2(REG2_REG_8__SCAN_IN),
.A1(n12357),
.ZN(n12358));
NAND2_X1 U8303 (.A2(n12358),
.A1(n12359),
.ZN(n12360));
NAND2_X1 U8304 (.A2(REG2_REG_9__SCAN_IN),
.A1(n12360),
.ZN(n12116));
NAND3_X1 U8305 (.A3(n12397),
.A1(n13798),
.A2(n12398),
.ZN(n12361));
NAND2_X1 U8306 (.A2(n12361),
.A1(jexoRSiRmgnTTbxiBcsGLhbKTivhVojg_Z),
.ZN(n12368));
NAND2_X1 U8307 (.A2(n12392),
.A1(n12393),
.ZN(n12363));
NAND2_X1 U8308 (.A2(n13804),
.A1(n12363),
.ZN(n12366));
NAND2_X1 U8309 (.A2(n12397),
.A1(n12398),
.ZN(n12364));
NAND2_X1 U8310 (.A2(n12364),
.A1(n13798),
.ZN(n12365));
NAND3_X1 U8311 (.A3(n13801),
.A1(n12366),
.A2(n12365),
.ZN(n12367));
MUX2_X1 U8312 (.S(n13773),
.A(n12368),
.B(n12367),
.Z(n12369));
AOI211_X1 U8313 (.C1(FE_OFN1_n13320),
.A(n12370),
.C2(ADDR_REG_9__SCAN_IN),
.B(n12369),
.ZN(n12371));
INV_X1 U8314 (.A(n12371),
.ZN(U3249));
INV_X1 U8316 (.A(n12374),
.ZN(n12373));
MUX2_X1 U8317 (.S(n12372),
.A(n12374),
.B(n12373),
.Z(n12383));
XNOR2_X1 U8318 (.B(n12375),
.A(n12379),
.ZN(n12376));
XNOR2_X1 U8319 (.B(n12376),
.A(n12377),
.ZN(n12381));
NAND2_X1 U8320 (.A2(ADDR_REG_7__SCAN_IN),
.A1(FE_OFN1_n13320),
.ZN(n12378));
NAND2_X1 U8321 (.A2(REG3_REG_7__SCAN_IN),
.A1(U3149),
.ZN(n12651));
OAI211_X1 U8322 (.C1(n13801),
.A(n12378),
.C2(n12379),
.B(n12651),
.ZN(n12380));
AOI21_X1 U8323 (.A(n12380),
.B2(n12381),
.B1(n13798),
.ZN(n12382));
OAI21_X1 U8324 (.A(n12382),
.B2(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.B1(n12383),
.ZN(U3247));
INV_X1 U8325 (.A(n12384),
.ZN(n12385));
NOR2_X1 U8326 (.A2(n12385),
.A1(n12386),
.ZN(n12388));
XNOR2_X1 U8327 (.B(n12387),
.A(n12388),
.ZN(n12391));
AOI22_X1 U8328 (.B2(n13784),
.B1(n13035),
.A1(n13038),
.A2(n11358),
.ZN(n12390));
AOI22_X1 U8329 (.B2(n13132),
.B1(n13037),
.A1(n12860),
.A2(REG3_REG_2__SCAN_IN),
.ZN(n12389));
OAI211_X1 U8330 (.C1(n12391),
.A(n12390),
.C2(n13005),
.B(n12389),
.ZN(U3234));
AND2_X1 U8331 (.A2(REG3_REG_11__SCAN_IN),
.A1(U3149),
.ZN(n12604));
NAND2_X1 U8332 (.A2(n13773),
.A1(n12392),
.ZN(n12394));
NAND2_X1 U8333 (.A2(n12393),
.A1(n12394),
.ZN(n13239));
OR2_X1 U8334 (.A2(REG1_REG_10__SCAN_IN),
.A1(n13772),
.ZN(n12395));
NAND2_X1 U8336 (.A2(n12396),
.A1(n12397),
.ZN(n12399));
NAND2_X1 U8337 (.A2(n12398),
.A1(n12399),
.ZN(n13240));
NOR2_X1 U8338 (.A2(REG2_REG_10__SCAN_IN),
.A1(n13772),
.ZN(n12400));
XNOR2_X1 U8341 (.B(REG2_REG_11__SCAN_IN),
.A(n12584),
.ZN(n12404));
OAI22_X1 U8342 (.B2(n13795),
.B1(n12404),
.A1(n12403),
.A2(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.ZN(n12408));
INV_X1 U8343 (.A(n12403),
.ZN(n12406));
AOI21_X1 U8345 (.A(n13292),
.B2(n13798),
.B1(n12404),
.ZN(n12405));
OAI21_X1 U8346 (.A(n12405),
.B2(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.B1(n12406),
.ZN(n12407));
MUX2_X1 U8347 (.S(n13771),
.A(n12408),
.B(n12407),
.Z(n12409));
AOI211_X1 U8348 (.C1(FE_OFN1_n13320),
.A(n12604),
.C2(ADDR_REG_11__SCAN_IN),
.B(n12409),
.ZN(n12410));
INV_X1 U8349 (.A(n12410),
.ZN(U3251));
OAI22_X1 U8350 (.B2(n12413),
.B1(STATE_REG_SCAN_IN),
.A1(n12990),
.A2(n13131),
.ZN(n12414));
INV_X1 U8351 (.A(n12414),
.ZN(n12416));
AOI22_X1 U8352 (.B2(n12490),
.B1(n13037),
.A1(n13035),
.A2(n13221),
.ZN(n12415));
OAI211_X1 U8353 (.C1(n13041),
.A(n12416),
.C2(REG3_REG_3__SCAN_IN),
.B(n12415),
.ZN(n12417));
AOI21_X1 U8354 (.A(n12417),
.B2(n13043),
.B1(n12418),
.ZN(n12419));
INV_X1 U8355 (.A(n12419),
.ZN(U3215));
INV_X1 U8356 (.A(n12421),
.ZN(n12422));
XNOR2_X1 U8357 (.B(n12422),
.A(n12420),
.ZN(n12516));
OAI22_X1 U8358 (.B2(n13698),
.B1(n12423),
.A1(n13819),
.A2(n12424),
.ZN(n12427));
XNOR2_X1 U8359 (.B(n13122),
.A(n12420),
.ZN(n12425));
AOI22_X1 U8360 (.B2(FE_OFN20_n11698),
.B1(n13690),
.A1(n12425),
.A2(n13672),
.ZN(n12518));
INV_X1 U8361 (.A(n12518),
.ZN(n12426));
AOI211_X1 U8362 (.C1(n13829),
.A(n12427),
.C2(n12516),
.B(n12426),
.ZN(n12489));
INV_X1 U8363 (.A(FE_OFN7_n13835),
.ZN(n13649));
INV_X1 U8364 (.A(n12428),
.ZN(n12431));
NAND2_X1 U8365 (.A2(n12429),
.A1(n11842),
.ZN(n12430));
NAND2_X1 U8366 (.A2(n12430),
.A1(n12431),
.ZN(n12514));
INV_X1 U8367 (.A(n12514),
.ZN(n12487));
AOI22_X1 U8368 (.B2(REG1_REG_1__SCAN_IN),
.B1(n13839),
.A1(n13649),
.A2(n12487),
.ZN(n12432));
OAI21_X1 U8369 (.A(n12432),
.B2(n13839),
.B1(n12489),
.ZN(U3519));
XNOR2_X1 U8370 (.B(n12434),
.A(n12433),
.ZN(n12493));
INV_X1 U8371 (.A(n12434),
.ZN(n13097));
XNOR2_X1 U8372 (.B(n13097),
.A(n12435),
.ZN(n12436));
AOI22_X1 U8373 (.B2(n13221),
.B1(n13690),
.A1(n12436),
.A2(n13672),
.ZN(n12497));
AOI22_X1 U8374 (.B2(n12490),
.B1(n13623),
.A1(n13688),
.A2(FE_OFN20_n11698),
.ZN(n12437));
OAI211_X1 U8375 (.C1(n13619),
.A(n12497),
.C2(n12493),
.B(n12437),
.ZN(n12701));
INV_X1 U8378 (.A(n12496),
.ZN(n12699));
OAI22_X1 U8379 (.B2(n12441),
.B1(n13841),
.A1(FE_OFN7_n13835),
.A2(n12699),
.ZN(n12442));
AOI21_X1 U8380 (.A(n12442),
.B2(n13841),
.B1(n12701),
.ZN(n12443));
INV_X1 U8381 (.A(n12443),
.ZN(U3521));
INV_X1 U8384 (.A(n12451),
.ZN(n13845));
XNOR2_X1 U8385 (.B(n13083),
.A(n12446),
.ZN(n12449));
AOI22_X1 U8386 (.B2(n13784),
.B1(n13690),
.A1(n13688),
.A2(n11358),
.ZN(n12448));
NAND2_X1 U8387 (.A2(n13132),
.A1(n13623),
.ZN(n12447));
OAI211_X1 U8388 (.C1(n12449),
.A(n12448),
.C2(n13568),
.B(n12447),
.ZN(n12450));
AOI21_X1 U8389 (.A(n12450),
.B2(n12451),
.B1(n12452),
.ZN(n13850));
OAI21_X1 U8390 (.A(n13850),
.B2(n13845),
.B1(n12453),
.ZN(n12705));
OAI21_X1 U8391 (.A(n12439),
.B2(n13128),
.B1(n12428),
.ZN(n13843));
OAI22_X1 U8392 (.B2(n12454),
.B1(n13841),
.A1(FE_OFN7_n13835),
.A2(n13843),
.ZN(n12455));
AOI21_X1 U8393 (.A(n12455),
.B2(n13841),
.B1(n12705),
.ZN(n12456));
INV_X1 U8394 (.A(n12456),
.ZN(U3520));
XNOR2_X1 U8395 (.B(n13138),
.A(n13818),
.ZN(n13084));
XNOR2_X1 U8396 (.B(n13084),
.A(n12457),
.ZN(n12458));
AOI222_X1 U8397 (.C2(n13690),
.C1(n13220),
.B2(n13623),
.B1(n13138),
.A1(n13672),
.A2(n12458),
.ZN(n13792));
XOR2_X1 U8398 (.B(n13084),
.A(n12459),
.Z(n13790));
AOI22_X1 U8399 (.B2(n13784),
.B1(n13688),
.A1(n13790),
.A2(n13829),
.ZN(n12460));
NAND2_X1 U8400 (.A2(n12460),
.A1(n13792),
.ZN(n12730));
OR2_X1 U8401 (.A2(n13135),
.A1(n12438),
.ZN(n12462));
NAND2_X1 U8402 (.A2(n12462),
.A1(n12461),
.ZN(n13787));
OAI22_X1 U8403 (.B2(n12463),
.B1(n13841),
.A1(FE_OFN7_n13835),
.A2(n13787),
.ZN(n12464));
AOI21_X1 U8404 (.A(n12464),
.B2(n13841),
.B1(n12730),
.ZN(n12465));
INV_X1 U8405 (.A(n12465),
.ZN(U3522));
NAND2_X1 U8406 (.A2(n12466),
.A1(n12536),
.ZN(n12467));
XNOR2_X1 U8407 (.B(n12467),
.A(n12614),
.ZN(n12472));
AOI21_X1 U8408 (.A(n12468),
.B2(n13784),
.B1(n13038),
.ZN(n12470));
AOI22_X1 U8409 (.B2(n13138),
.B1(n13037),
.A1(n13035),
.A2(n13220),
.ZN(n12469));
OAI211_X1 U8410 (.C1(n13041),
.A(n12470),
.C2(n13780),
.B(n12469),
.ZN(n12471));
AOI21_X1 U8411 (.A(n12471),
.B2(n13043),
.B1(n12472),
.ZN(n12473));
INV_X1 U8412 (.A(n12473),
.ZN(U3227));
XNOR2_X1 U8413 (.B(n12474),
.A(n13094),
.ZN(n12475));
OAI222_X1 U8414 (.C2(n12652),
.C1(n13627),
.B2(n13568),
.B1(n12475),
.A1(n13698),
.A2(n11795),
.ZN(n13820));
INV_X1 U8415 (.A(n13820),
.ZN(n12486));
INV_X1 U8416 (.A(n12476),
.ZN(n12479));
AOI211_X1 U8417 (.C1(n12459),
.A(n12477),
.C2(n13084),
.B(n13094),
.ZN(n12478));
NOR2_X1 U8418 (.A2(n12478),
.A1(n12479),
.ZN(n13822));
NAND2_X1 U8419 (.A2(n12543),
.A1(n12461),
.ZN(n12481));
NAND2_X1 U8420 (.A2(n12481),
.A1(n12480),
.ZN(n13834));
OAI22_X1 U8421 (.B2(n13779),
.B1(n12546),
.A1(n13782),
.A2(n11395),
.ZN(n12482));
AOI21_X1 U8422 (.A(n12482),
.B2(n13221),
.B1(n13785),
.ZN(n12483));
OAI21_X1 U8423 (.A(n12483),
.B2(n13834),
.B1(n13844),
.ZN(n12484));
AOI21_X1 U8424 (.A(n12484),
.B2(n13789),
.B1(n13822),
.ZN(n12485));
OAI21_X1 U8425 (.A(n12485),
.B2(n11157),
.B1(n12486),
.ZN(U3285));
AOI22_X1 U8426 (.B2(REG0_REG_1__SCAN_IN),
.B1(n13860),
.A1(n13729),
.A2(n12487),
.ZN(n12488));
OAI21_X1 U8427 (.A(n12488),
.B2(n13860),
.B1(n12489),
.ZN(U3469));
NAND2_X1 U8428 (.A2(FE_OFN20_n11698),
.A1(n13785),
.ZN(n12492));
NAND2_X1 U8429 (.A2(n12490),
.A1(FE_OFN8_n11821),
.ZN(n12491));
OAI211_X1 U8430 (.C1(n13779),
.A(n12492),
.C2(REG3_REG_3__SCAN_IN),
.B(n12491),
.ZN(n12495));
NOR2_X1 U8431 (.A2(n12493),
.A1(n13584),
.ZN(n12494));
AOI211_X1 U8432 (.C1(FE_OFN2_n13580),
.A(n12495),
.C2(n12496),
.B(n12494),
.ZN(n12500));
MUX2_X1 U8433 (.S(n13782),
.A(n12498),
.B(n12497),
.Z(n12499));
NAND2_X1 U8434 (.A2(n12499),
.A1(n12500),
.ZN(U3287));
INV_X1 U8435 (.A(n13374),
.ZN(n12502));
AOI211_X1 U8436 (.C1(n12620),
.A(n12502),
.C2(n12480),
.B(n11295),
.ZN(n13828));
NAND2_X1 U8437 (.A2(n13139),
.A1(n13086),
.ZN(n12507));
XOR2_X1 U8438 (.B(n12523),
.A(n12507),
.Z(n12505));
OAI22_X1 U8439 (.B2(n12618),
.B1(n13819),
.A1(n12675),
.A2(n13627),
.ZN(n12503));
AOI21_X1 U8440 (.A(n12503),
.B2(n13623),
.B1(n12620),
.ZN(n12504));
OAI21_X1 U8441 (.A(n12504),
.B2(n13568),
.B1(n12505),
.ZN(n13827));
AOI21_X1 U8442 (.A(n13827),
.B2(n13315),
.B1(n13828),
.ZN(n12511));
INV_X1 U8443 (.A(n12506),
.ZN(n12521));
XNOR2_X1 U8444 (.B(n12507),
.A(n12521),
.ZN(n13830));
OAI22_X1 U8445 (.B2(n13779),
.B1(n12623),
.A1(n13782),
.A2(n12508),
.ZN(n12509));
AOI21_X1 U8446 (.A(n12509),
.B2(n13789),
.B1(n13830),
.ZN(n12510));
OAI21_X1 U8447 (.A(n12510),
.B2(n11157),
.B1(n12511),
.ZN(U3284));
AOI22_X1 U8448 (.B2(n11831),
.B1(n13785),
.A1(n11842),
.A2(FE_OFN8_n11821),
.ZN(n12513));
AOI22_X1 U8449 (.B2(REG3_REG_1__SCAN_IN),
.B1(n13842),
.A1(n11157),
.A2(REG2_REG_1__SCAN_IN),
.ZN(n12512));
OAI211_X1 U8450 (.C1(n13844),
.A(n12513),
.C2(n12514),
.B(n12512),
.ZN(n12515));
AOI21_X1 U8451 (.A(n12515),
.B2(n12516),
.B1(n13789),
.ZN(n12517));
OAI21_X1 U8452 (.A(n12517),
.B2(n12518),
.B1(n11157),
.ZN(U3289));
AOI21_X1 U8453 (.A(n12620),
.B2(n13219),
.B1(n12506),
.ZN(n12520));
AOI21_X1 U8454 (.A(n12520),
.B2(n12521),
.B1(n12652),
.ZN(n12522));
XNOR2_X1 U8455 (.B(n12522),
.A(n12526),
.ZN(n12639));
NAND2_X1 U8456 (.A2(n13086),
.A1(n12523),
.ZN(n12524));
NAND2_X1 U8457 (.A2(n13139),
.A1(n12524),
.ZN(n12525));
XNOR2_X1 U8458 (.B(n12525),
.A(n12526),
.ZN(n12641));
NAND2_X1 U8459 (.A2(FE_OFN9_n13503),
.A1(n12641),
.ZN(n12534));
XNOR2_X1 U8460 (.B(n12654),
.A(n12501),
.ZN(n12724));
INV_X1 U8461 (.A(n12724),
.ZN(n12532));
AOI22_X1 U8462 (.B2(n13217),
.B1(FE_OFN10_n13571),
.A1(FE_OFN8_n11821),
.A2(n12654),
.ZN(n12530));
INV_X1 U8463 (.A(n12657),
.ZN(n12528));
AOI22_X1 U8464 (.B2(n12528),
.B1(n13842),
.A1(n11157),
.A2(REG2_REG_7__SCAN_IN),
.ZN(n12529));
OAI211_X1 U8465 (.C1(n12652),
.A(n12530),
.C2(n13577),
.B(n12529),
.ZN(n12531));
AOI21_X1 U8466 (.A(n12531),
.B2(n12532),
.B1(FE_OFN2_n13580),
.ZN(n12533));
OAI211_X1 U8467 (.C1(n13584),
.A(n12534),
.C2(n12639),
.B(n12533),
.ZN(U3283));
AOI21_X1 U8468 (.A(n12535),
.B2(n12536),
.B1(n12614),
.ZN(n12540));
NAND2_X1 U8469 (.A2(n12537),
.A1(n12538),
.ZN(n12539));
XOR2_X1 U8470 (.B(n12539),
.A(n12540),
.Z(n12548));
OAI21_X1 U8471 (.A(n12541),
.B2(n13818),
.B1(n12990),
.ZN(n12542));
INV_X1 U8472 (.A(n12542),
.ZN(n12545));
AOI22_X1 U8473 (.B2(n12543),
.B1(n13037),
.A1(n13035),
.A2(n13219),
.ZN(n12544));
OAI211_X1 U8474 (.C1(n13041),
.A(n12545),
.C2(n12546),
.B(n12544),
.ZN(n12547));
AOI21_X1 U8475 (.A(n12547),
.B2(n13043),
.B1(n12548),
.ZN(n12549));
INV_X1 U8476 (.A(n12549),
.ZN(U3224));
NOR2_X1 U8477 (.A2(FE_OFN9_n13503),
.A1(n13789),
.ZN(n12555));
OAI22_X1 U8478 (.B2(n13779),
.B1(n12550),
.A1(n13782),
.A2(n12551),
.ZN(n12553));
AOI21_X1 U8479 (.A(n12863),
.B2(n13844),
.B1(n13518),
.ZN(n12552));
AOI211_X1 U8480 (.C1(FE_OFN10_n13571),
.A(n12553),
.C2(n11358),
.B(n12552),
.ZN(n12554));
OAI21_X1 U8481 (.A(n12554),
.B2(n12555),
.B1(n13078),
.ZN(U3290));
OAI21_X1 U8490 (.A(n12563),
.B2(n12629),
.B1(n12564),
.ZN(n12698));
AOI22_X1 U8491 (.B2(n11157),
.B1(REG2_REG_8__SCAN_IN),
.A1(FE_OFN8_n11821),
.A2(n12677),
.ZN(n12566));
AOI22_X1 U8492 (.B2(n13216),
.B1(FE_OFN10_n13571),
.A1(n13785),
.A2(n13218),
.ZN(n12565));
OAI211_X1 U8493 (.C1(n12698),
.A(n12566),
.C2(n13844),
.B(n12565),
.ZN(n12567));
AOI21_X1 U8494 (.A(n12567),
.B2(n13789),
.B1(n12631),
.ZN(n12568));
OAI21_X1 U8495 (.A(n12568),
.B2(n11157),
.B1(n12569),
.ZN(U3282));
NAND2_X1 U8497 (.A2(n13771),
.A1(n12570),
.ZN(n12574));
INV_X1 U8498 (.A(n12571),
.ZN(n12572));
NAND2_X1 U8499 (.A2(REG1_REG_11__SCAN_IN),
.A1(n12572),
.ZN(n12573));
NAND2_X1 U8500 (.A2(n12573),
.A1(n12574),
.ZN(n13250));
NAND2_X1 U8501 (.A2(REG1_REG_12__SCAN_IN),
.A1(n13250),
.ZN(n12576));
NAND2_X1 U8502 (.A2(n12576),
.A1(n12577),
.ZN(n13263));
INV_X1 U8503 (.A(n13269),
.ZN(n12578));
OAI21_X1 U8504 (.A(n12578),
.B2(REG1_REG_13__SCAN_IN),
.B1(n13263),
.ZN(n12580));
NAND2_X1 U8505 (.A2(REG1_REG_13__SCAN_IN),
.A1(n13263),
.ZN(n12579));
OR2_X1 U8506 (.A2(REG1_REG_14__SCAN_IN),
.A1(n13770),
.ZN(n12581));
XNOR2_X1 U8508 (.B(n12773),
.A(n12582),
.ZN(n12599));
NAND2_X1 U8511 (.A2(REG2_REG_11__SCAN_IN),
.A1(n13771),
.ZN(n12585));
NAND2_X1 U8512 (.A2(n12585),
.A1(n12586),
.ZN(n12587));
NAND2_X1 U8513 (.A2(REG2_REG_12__SCAN_IN),
.A1(n12587),
.ZN(n13254));
NAND2_X1 U8514 (.A2(n13257),
.A1(n13254),
.ZN(n12588));
NAND2_X1 U8515 (.A2(n13253),
.A1(n12588),
.ZN(n13264));
AND2_X1 U8516 (.A2(n12589),
.A1(n13269),
.ZN(n12590));
NAND2_X1 U8520 (.A2(REG2_REG_14__SCAN_IN),
.A1(n13770),
.ZN(n12592));
NAND2_X1 U8521 (.A2(n12592),
.A1(n12593),
.ZN(n12765));
XNOR2_X1 U8522 (.B(REG2_REG_15__SCAN_IN),
.A(n12766),
.ZN(n12594));
XNOR2_X1 U8523 (.B(n12594),
.A(n12765),
.ZN(n12597));
AND2_X1 U8524 (.A2(REG3_REG_15__SCAN_IN),
.A1(U3149),
.ZN(n13034));
AOI21_X1 U8525 (.A(n13034),
.B2(ADDR_REG_15__SCAN_IN),
.B1(FE_OFN1_n13320),
.ZN(n12595));
OAI21_X1 U8526 (.A(n12595),
.B2(n13801),
.B1(n12773),
.ZN(n12596));
AOI21_X1 U8527 (.A(n12596),
.B2(n13798),
.B1(n12597),
.ZN(n12598));
OAI21_X1 U8528 (.A(n12598),
.B2(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.B1(n12599),
.ZN(U3255));
XNOR2_X1 U8530 (.B(n12600),
.A(n12603),
.ZN(n12608));
AOI21_X1 U8531 (.A(n12604),
.B2(n13214),
.B1(n13035),
.ZN(n12606));
AOI22_X1 U8532 (.B2(n12822),
.B1(n13037),
.A1(n13038),
.A2(n13215),
.ZN(n12605));
OAI211_X1 U8533 (.C1(n13041),
.A(n12606),
.C2(n12818),
.B(n12605),
.ZN(n12607));
AOI21_X1 U8534 (.A(n12607),
.B2(n13043),
.B1(n12608),
.ZN(n12609));
INV_X1 U8535 (.A(n12609),
.ZN(U3233));
INV_X1 U8536 (.A(n12610),
.ZN(n12613));
INV_X1 U8537 (.A(n12611),
.ZN(n12612));
AOI21_X1 U8538 (.A(n12612),
.B2(n12613),
.B1(n12614),
.ZN(n12646));
NAND2_X1 U8539 (.A2(n12644),
.A1(n12615),
.ZN(n12616));
XOR2_X1 U8540 (.B(n12616),
.A(n12646),
.Z(n12625));
OAI21_X1 U8541 (.A(n12617),
.B2(n12618),
.B1(n12990),
.ZN(n12619));
INV_X1 U8542 (.A(n12619),
.ZN(n12622));
AOI22_X1 U8543 (.B2(n12620),
.B1(n13037),
.A1(n13035),
.A2(n13218),
.ZN(n12621));
OAI211_X1 U8544 (.C1(n13041),
.A(n12622),
.C2(n12623),
.B(n12621),
.ZN(n12624));
AOI21_X1 U8545 (.A(n12624),
.B2(n13043),
.B1(n12625),
.ZN(n12626));
INV_X1 U8546 (.A(n12626),
.ZN(U3236));
NAND2_X1 U8547 (.A2(n13218),
.A1(n13688),
.ZN(n12628));
NAND2_X1 U8548 (.A2(n13216),
.A1(n13690),
.ZN(n12627));
OAI211_X1 U8549 (.C1(n13698),
.A(n12628),
.C2(n12629),
.B(n12627),
.ZN(n12630));
AOI21_X1 U8550 (.A(n12630),
.B2(n13829),
.B1(n12631),
.ZN(n12632));
NAND2_X1 U8551 (.A2(n12632),
.A1(n12633),
.ZN(n12695));
INV_X1 U8552 (.A(n12695),
.ZN(n12634));
MUX2_X1 U8553 (.S(FE_OFN3_n13832),
.A(n12635),
.B(n12634),
.Z(n12636));
OAI21_X1 U8554 (.A(n12636),
.B2(FE_OFN21_n13759),
.B1(n12698),
.ZN(U3483));
OAI22_X1 U8555 (.B2(n12828),
.B1(n13627),
.A1(n12652),
.A2(n13819),
.ZN(n12637));
AOI21_X1 U8556 (.A(n12637),
.B2(n13623),
.B1(n12654),
.ZN(n12638));
OAI21_X1 U8557 (.A(n12638),
.B2(n13619),
.B1(n12639),
.ZN(n12640));
AOI21_X1 U8558 (.A(n12640),
.B2(n12641),
.B1(n13672),
.ZN(n12727));
MUX2_X1 U8559 (.S(n13841),
.A(n12642),
.B(n12727),
.Z(n12643));
OAI21_X1 U8560 (.A(n12643),
.B2(FE_OFN7_n13835),
.B1(n12724),
.ZN(U3525));
OAI21_X1 U8561 (.A(n12644),
.B2(n12645),
.B1(n12646),
.ZN(n12650));
NAND2_X1 U8562 (.A2(n12647),
.A1(n12648),
.ZN(n12649));
XNOR2_X1 U8563 (.B(n12649),
.A(n12650),
.ZN(n12659));
OAI21_X1 U8564 (.A(n12651),
.B2(n12652),
.B1(n12990),
.ZN(n12653));
INV_X1 U8565 (.A(n12653),
.ZN(n12656));
AOI22_X1 U8566 (.B2(n12654),
.B1(n13037),
.A1(n13035),
.A2(n13217),
.ZN(n12655));
OAI211_X1 U8567 (.C1(n13041),
.A(n12656),
.C2(n12657),
.B(n12655),
.ZN(n12658));
AOI21_X1 U8568 (.A(n12658),
.B2(n13043),
.B1(n12659),
.ZN(n12660));
INV_X1 U8569 (.A(n12660),
.ZN(U3210));
AND2_X1 U8570 (.A2(REG3_REG_14__SCAN_IN),
.A1(U3149),
.ZN(n12900));
XNOR2_X1 U8571 (.B(REG1_REG_14__SCAN_IN),
.A(n12661),
.ZN(n12663));
XNOR2_X1 U8572 (.B(REG2_REG_14__SCAN_IN),
.A(n12662),
.ZN(n12664));
OAI22_X1 U8573 (.B2(n13795),
.B1(n12664),
.A1(n12663),
.A2(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.ZN(n12668));
INV_X1 U8574 (.A(n12663),
.ZN(n12666));
AOI21_X1 U8575 (.A(n13292),
.B2(n13798),
.B1(n12664),
.ZN(n12665));
OAI21_X1 U8576 (.A(n12665),
.B2(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.B1(n12666),
.ZN(n12667));
MUX2_X1 U8577 (.S(n13770),
.A(n12668),
.B(n12667),
.Z(n12669));
AOI211_X1 U8578 (.C1(FE_OFN1_n13320),
.A(n12900),
.C2(ADDR_REG_14__SCAN_IN),
.B(n12669),
.ZN(n12670));
INV_X1 U8579 (.A(n12670),
.ZN(U3254));
INV_X1 U8580 (.A(n12671),
.ZN(n12750));
NAND2_X1 U8581 (.A2(n12672),
.A1(n12749),
.ZN(n12673));
XNOR2_X1 U8582 (.B(n12673),
.A(n12750),
.ZN(n12682));
OAI21_X1 U8583 (.A(n12674),
.B2(n12675),
.B1(n12990),
.ZN(n12676));
INV_X1 U8584 (.A(n12676),
.ZN(n12679));
AOI22_X1 U8585 (.B2(n12677),
.B1(n13037),
.A1(n13035),
.A2(n13216),
.ZN(n12678));
OAI211_X1 U8586 (.C1(n13041),
.A(n12679),
.C2(n12680),
.B(n12678),
.ZN(n12681));
AOI21_X1 U8587 (.A(n12681),
.B2(n13043),
.B1(n12682),
.ZN(n12683));
INV_X1 U8588 (.A(n12683),
.ZN(U3218));
NAND2_X1 U8589 (.A2(n13150),
.A1(n11173),
.ZN(n13088));
XOR2_X1 U8590 (.B(n13088),
.A(n12684),
.Z(n12685));
OAI22_X1 U8591 (.B2(n13627),
.B1(n13700),
.A1(n12685),
.A2(n13568),
.ZN(n12829));
INV_X1 U8592 (.A(n12829),
.ZN(n12694));
XNOR2_X1 U8593 (.B(n13088),
.A(n12686),
.ZN(n12831));
NAND2_X1 U8594 (.A2(n12757),
.A1(n12563),
.ZN(n12687));
NAND2_X1 U8595 (.A2(n12687),
.A1(n12712),
.ZN(n12837));
INV_X1 U8596 (.A(n12760),
.ZN(n12688));
AOI22_X1 U8597 (.B2(n12688),
.B1(n13842),
.A1(n11157),
.A2(REG2_REG_9__SCAN_IN),
.ZN(n12689));
OAI21_X1 U8598 (.A(n12689),
.B2(n12828),
.B1(n13577),
.ZN(n12690));
AOI21_X1 U8599 (.A(n12690),
.B2(FE_OFN8_n11821),
.B1(n12757),
.ZN(n12691));
OAI21_X1 U8600 (.A(n12691),
.B2(n13844),
.B1(n12837),
.ZN(n12692));
AOI21_X1 U8601 (.A(n12692),
.B2(n13789),
.B1(n12831),
.ZN(n12693));
OAI21_X1 U8602 (.A(n12693),
.B2(n11157),
.B1(n12694),
.ZN(U3281));
MUX2_X1 U8603 (.S(n13839),
.A(n12695),
.B(REG1_REG_8__SCAN_IN),
.Z(n12696));
INV_X1 U8604 (.A(n12696),
.ZN(n12697));
OAI21_X1 U8605 (.A(n12697),
.B2(n12698),
.B1(FE_OFN7_n13835),
.ZN(U3526));
OAI22_X1 U8606 (.B2(n11376),
.B1(FE_OFN3_n13832),
.A1(FE_OFN21_n13759),
.A2(n12699),
.ZN(n12700));
AOI21_X1 U8607 (.A(n12700),
.B2(FE_OFN3_n13832),
.B1(n12701),
.ZN(n12702));
INV_X1 U8608 (.A(n12702),
.ZN(U3473));
OAI22_X1 U8609 (.B2(n12703),
.B1(FE_OFN3_n13832),
.A1(FE_OFN21_n13759),
.A2(n13843),
.ZN(n12704));
AOI21_X1 U8610 (.A(n12704),
.B2(FE_OFN3_n13832),
.B1(n12705),
.ZN(n12706));
INV_X1 U8611 (.A(n12706),
.ZN(U3471));
NAND2_X1 U8612 (.A2(n12707),
.A1(n12686),
.ZN(n12709));
NAND2_X1 U8613 (.A2(n12708),
.A1(n12709),
.ZN(n12710));
XNOR2_X1 U8614 (.B(n13098),
.A(n12710),
.ZN(n12798));
XNOR2_X1 U8615 (.B(n13098),
.A(n12711),
.ZN(n12800));
NAND2_X1 U8616 (.A2(FE_OFN9_n13503),
.A1(n12800),
.ZN(n12722));
INV_X1 U8617 (.A(n12713),
.ZN(n12714));
OAI21_X1 U8618 (.A(n12714),
.B2(n12718),
.B1(n11192),
.ZN(n12806));
INV_X1 U8619 (.A(n12806),
.ZN(n12720));
AOI22_X1 U8620 (.B2(n13687),
.B1(FE_OFN10_n13571),
.A1(n13785),
.A2(n13216),
.ZN(n12717));
INV_X1 U8621 (.A(n12744),
.ZN(n12715));
AOI22_X1 U8622 (.B2(n12715),
.B1(n13842),
.A1(n11157),
.A2(REG2_REG_10__SCAN_IN),
.ZN(n12716));
OAI211_X1 U8623 (.C1(n12718),
.A(n12717),
.C2(n13518),
.B(n12716),
.ZN(n12719));
AOI21_X1 U8624 (.A(n12719),
.B2(FE_OFN2_n13580),
.B1(n12720),
.ZN(n12721));
OAI211_X1 U8625 (.C1(n13584),
.A(n12722),
.C2(n12798),
.B(n12721),
.ZN(U3280));
INV_X1 U8626 (.A(REG0_REG_7__SCAN_IN),
.ZN(n12723));
OAI22_X1 U8627 (.B2(n12723),
.B1(FE_OFN3_n13832),
.A1(n12724),
.A2(FE_OFN21_n13759),
.ZN(n12725));
INV_X1 U8628 (.A(n12725),
.ZN(n12726));
OAI21_X1 U8629 (.A(n12726),
.B2(n13860),
.B1(n12727),
.ZN(U3481));
OAI22_X1 U8630 (.B2(n12728),
.B1(FE_OFN3_n13832),
.A1(FE_OFN21_n13759),
.A2(n13787),
.ZN(n12729));
AOI21_X1 U8631 (.A(n12729),
.B2(FE_OFN3_n13832),
.B1(n12730),
.ZN(n12731));
INV_X1 U8632 (.A(n12731),
.ZN(U3475));
INV_X1 U8633 (.A(n12732),
.ZN(n12735));
INV_X1 U8634 (.A(n12733),
.ZN(n12734));
AOI21_X1 U8635 (.A(n12734),
.B2(n12735),
.B1(n12750),
.ZN(n12740));
INV_X1 U8636 (.A(n12736),
.ZN(n12738));
NAND2_X1 U8637 (.A2(n12737),
.A1(n12738),
.ZN(n12739));
XOR2_X1 U8638 (.B(n12739),
.A(n12740),
.Z(n12746));
NAND2_X1 U8639 (.A2(REG3_REG_10__SCAN_IN),
.A1(U3149),
.ZN(n13248));
OAI21_X1 U8640 (.A(n13248),
.B2(n12794),
.B1(n12990),
.ZN(n12741));
INV_X1 U8641 (.A(n12741),
.ZN(n12743));
AOI22_X1 U8642 (.B2(n12796),
.B1(n13037),
.A1(n13035),
.A2(n13687),
.ZN(n12742));
OAI211_X1 U8643 (.C1(n13041),
.A(n12743),
.C2(n12744),
.B(n12742),
.ZN(n12745));
AOI21_X1 U8644 (.A(n12745),
.B2(n13043),
.B1(n12746),
.ZN(n12747));
INV_X1 U8645 (.A(n12747),
.ZN(U3214));
AOI21_X1 U8646 (.A(n12748),
.B2(n12749),
.B1(n12750),
.ZN(n12754));
NAND2_X1 U8647 (.A2(n12751),
.A1(n12752),
.ZN(n12753));
XOR2_X1 U8648 (.B(n12753),
.A(n12754),
.Z(n12762));
OAI21_X1 U8649 (.A(n12755),
.B2(n12828),
.B1(n12990),
.ZN(n12756));
INV_X1 U8650 (.A(n12756),
.ZN(n12759));
AOI22_X1 U8651 (.B2(n12757),
.B1(n13037),
.A1(n13035),
.A2(n13215),
.ZN(n12758));
OAI211_X1 U8652 (.C1(n13041),
.A(n12759),
.C2(n12760),
.B(n12758),
.ZN(n12761));
AOI21_X1 U8653 (.A(n12761),
.B2(n13043),
.B1(n12762),
.ZN(n12763));
INV_X1 U8654 (.A(n12763),
.ZN(U3228));
INV_X1 U8657 (.A(n12770),
.ZN(n12769));
OR2_X1 U8658 (.A2(REG2_REG_15__SCAN_IN),
.A1(n12766),
.ZN(n12764));
NAND2_X1 U8659 (.A2(n12764),
.A1(n12765),
.ZN(n12768));
NAND2_X1 U8660 (.A2(REG2_REG_15__SCAN_IN),
.A1(n12766),
.ZN(n12767));
NAND2_X1 U8661 (.A2(n12767),
.A1(n12768),
.ZN(n13279));
MUX2_X1 U8662 (.S(n13279),
.A(n12770),
.B(n12769),
.Z(n12783));
INV_X1 U8663 (.A(REG1_REG_16__SCAN_IN),
.ZN(n13663));
XNOR2_X1 U8664 (.B(n13663),
.A(n13287),
.ZN(n12776));
AOI21_X1 U8665 (.A(n13292),
.B2(n13804),
.B1(n12776),
.ZN(n12779));
MUX2_X1 U8668 (.S(n13288),
.A(n12779),
.B(n12778),
.Z(n12782));
NAND2_X1 U8669 (.A2(REG3_REG_16__SCAN_IN),
.A1(U3149),
.ZN(n12963));
INV_X1 U8670 (.A(n12963),
.ZN(n12780));
AOI21_X1 U8671 (.A(n12780),
.B2(ADDR_REG_16__SCAN_IN),
.B1(FE_OFN1_n13320),
.ZN(n12781));
OAI211_X1 U8672 (.C1(n12783),
.A(n12782),
.C2(n13795),
.B(n12781),
.ZN(U3256));
XOR2_X1 U8673 (.B(n12784),
.A(n12785),
.Z(n12786));
XNOR2_X1 U8674 (.B(n12786),
.A(n12787),
.ZN(n12792));
NAND2_X1 U8675 (.A2(REG3_REG_12__SCAN_IN),
.A1(U3149),
.ZN(n13261));
OAI21_X1 U8676 (.A(n13261),
.B2(n13578),
.B1(n12990),
.ZN(n12788));
INV_X1 U8677 (.A(n12788),
.ZN(n12790));
AOI22_X1 U8678 (.B2(n13572),
.B1(n13037),
.A1(n13035),
.A2(n13689),
.ZN(n12789));
OAI211_X1 U8679 (.C1(n13041),
.A(n12790),
.C2(n13573),
.B(n12789),
.ZN(n12791));
AOI21_X1 U8680 (.A(n12791),
.B2(n13043),
.B1(n12792),
.ZN(n12793));
INV_X1 U8681 (.A(n12793),
.ZN(U3221));
INV_X1 U8682 (.A(REG0_REG_10__SCAN_IN),
.ZN(n12801));
OAI22_X1 U8683 (.B2(n13578),
.B1(n13627),
.A1(n12794),
.A2(n13819),
.ZN(n12795));
AOI21_X1 U8684 (.A(n12795),
.B2(n13623),
.B1(n12796),
.ZN(n12797));
OAI21_X1 U8685 (.A(n12797),
.B2(n13619),
.B1(n12798),
.ZN(n12799));
AOI21_X1 U8686 (.A(n12799),
.B2(n13672),
.B1(n12800),
.ZN(n12803));
MUX2_X1 U8687 (.S(FE_OFN3_n13832),
.A(n12801),
.B(n12803),
.Z(n12802));
OAI21_X1 U8688 (.A(n12802),
.B2(FE_OFN21_n13759),
.B1(n12806),
.ZN(U3487));
MUX2_X1 U8689 (.S(n13841),
.A(n12804),
.B(n12803),
.Z(n13737));
OAI21_X1 U8690 (.A(n12805),
.B2(n12806),
.B1(FE_OFN7_n13835),
.ZN(U3528));
XOR2_X1 U8691 (.B(n13095),
.A(n12808),
.Z(n12809));
OAI22_X1 U8692 (.B2(n13627),
.B1(n13680),
.A1(n12809),
.A2(n13568),
.ZN(n13701));
INV_X1 U8693 (.A(n13701),
.ZN(n12826));
NAND2_X1 U8694 (.A2(n12810),
.A1(n12686),
.ZN(n12813));
NAND2_X1 U8695 (.A2(n12811),
.A1(n12813),
.ZN(n12816));
AOI21_X1 U8697 (.A(n12815),
.B2(n12816),
.B1(n13095),
.ZN(n13703));
AND2_X1 U8698 (.A2(n13699),
.A1(n12713),
.ZN(n13570));
NOR2_X1 U8699 (.A2(n13699),
.A1(n12713),
.ZN(n12817));
INV_X1 U8700 (.A(REG2_REG_11__SCAN_IN),
.ZN(n12819));
OAI22_X1 U8701 (.B2(n13779),
.B1(n12818),
.A1(n13782),
.A2(n12819),
.ZN(n12821));
NOR2_X1 U8702 (.A2(n13700),
.A1(n13577),
.ZN(n12820));
AOI211_X1 U8703 (.C1(FE_OFN8_n11821),
.A(n12821),
.C2(n12822),
.B(n12820),
.ZN(n12823));
OAI21_X1 U8704 (.A(n12823),
.B2(n13844),
.B1(n13760),
.ZN(n12824));
AOI21_X1 U8705 (.A(n12824),
.B2(n13789),
.B1(n13703),
.ZN(n12825));
OAI21_X1 U8706 (.A(n12825),
.B2(n11157),
.B1(n12826),
.ZN(U3279));
OAI22_X1 U8707 (.B2(n13698),
.B1(n12827),
.A1(n13819),
.A2(n12828),
.ZN(n12830));
AOI211_X1 U8708 (.C1(n12831),
.A(n12830),
.C2(n13829),
.B(n12829),
.ZN(n12834));
MUX2_X1 U8709 (.S(FE_OFN3_n13832),
.A(n12832),
.B(n12834),
.Z(n12833));
OAI21_X1 U8710 (.A(n12833),
.B2(FE_OFN21_n13759),
.B1(n12837),
.ZN(U3485));
MUX2_X1 U8711 (.S(n13841),
.A(n12835),
.B(n12834),
.Z(n12836));
OAI21_X1 U8712 (.A(n12836),
.B2(n12837),
.B1(FE_OFN7_n13835),
.ZN(U3527));
INV_X1 U8713 (.A(IR_REG_30__SCAN_IN),
.ZN(n12838));
NAND2_X1 U8714 (.A2(n12838),
.A1(n12839),
.ZN(n12841));
INV_X1 U8715 (.A(DATAI_31_),
.ZN(n12840));
OAI22_X1 U8716 (.B2(n12840),
.B1(STATE_REG_SCAN_IN),
.A1(n11336),
.A2(n12841),
.ZN(U3321));
INV_X1 U8719 (.A(n12843),
.ZN(n12847));
INV_X1 U8720 (.A(REG2_REG_31__SCAN_IN),
.ZN(n12846));
NAND2_X1 U8721 (.A2(REG1_REG_31__SCAN_IN),
.A1(FE_DBTN1_n11467),
.ZN(n12845));
INV_X1 U8722 (.A(REG0_REG_31__SCAN_IN),
.ZN(n12868));
OR2_X1 U8723 (.A2(n12868),
.A1(n11418),
.ZN(n12844));
OAI211_X1 U8724 (.C1(n11469),
.A(n12845),
.C2(n12846),
.B(n12844),
.ZN(n13208));
NAND2_X1 U8725 (.A2(n13208),
.A1(n12847),
.ZN(n12867));
OAI21_X1 U8726 (.A(n12867),
.B2(n13698),
.B1(n12848),
.ZN(n12855));
NOR2_X1 U8727 (.A2(n12849),
.A1(FE_OFN3_n13832),
.ZN(n12850));
AOI21_X1 U8728 (.A(n12850),
.B2(n12855),
.B1(FE_OFN3_n13832),
.ZN(n12851));
OAI21_X1 U8729 (.A(n12851),
.B2(FE_OFN21_n13759),
.B1(n12858),
.ZN(U3516));
NOR2_X1 U8730 (.A2(n12852),
.A1(n13782),
.ZN(n12853));
AOI21_X1 U8731 (.A(n12853),
.B2(n12855),
.B1(n13782),
.ZN(n12854));
OAI21_X1 U8732 (.A(n12854),
.B2(n13844),
.B1(n12858),
.ZN(U3261));
NAND2_X1 U8733 (.A2(n12855),
.A1(n13841),
.ZN(n12857));
NAND2_X1 U8734 (.A2(REG1_REG_30__SCAN_IN),
.A1(n13839),
.ZN(n12856));
OAI211_X1 U8735 (.C1(n12858),
.A(n12857),
.C2(FE_OFN7_n13835),
.B(n12856),
.ZN(U3548));
NAND2_X1 U8736 (.A2(n13043),
.A1(n12859),
.ZN(n12862));
AOI22_X1 U8737 (.B2(n11358),
.B1(n13035),
.A1(REG3_REG_0__SCAN_IN),
.A2(n12860),
.ZN(n12861));
OAI211_X1 U8738 (.C1(n12991),
.A(n12862),
.C2(n12863),
.B(n12861),
.ZN(U3229));
NAND2_X1 U8739 (.A2(DATAI_31_),
.A1(n11569),
.ZN(n13069));
OAI21_X1 U8740 (.A(n12867),
.B2(n13698),
.B1(n13069),
.ZN(n12873));
NOR2_X1 U8741 (.A2(n12868),
.A1(FE_OFN3_n13832),
.ZN(n12869));
AOI21_X1 U8742 (.A(n12869),
.B2(n12873),
.B1(FE_OFN3_n13832),
.ZN(n12870));
OAI21_X1 U8743 (.A(n12870),
.B2(FE_OFN21_n13759),
.B1(n12876),
.ZN(U3517));
NAND2_X1 U8744 (.A2(n13782),
.A1(n12873),
.ZN(n12872));
NAND2_X1 U8745 (.A2(REG2_REG_31__SCAN_IN),
.A1(n11157),
.ZN(n12871));
OAI211_X1 U8746 (.C1(n12876),
.A(n12872),
.C2(n13844),
.B(n12871),
.ZN(U3260));
NAND2_X1 U8747 (.A2(n12873),
.A1(n13841),
.ZN(n12875));
NAND2_X1 U8748 (.A2(REG1_REG_31__SCAN_IN),
.A1(n13839),
.ZN(n12874));
OAI211_X1 U8749 (.C1(n12876),
.A(n12875),
.C2(FE_OFN7_n13835),
.B(n12874),
.ZN(U3549));
NAND2_X1 U8750 (.A2(n13785),
.A1(n13343),
.ZN(n12879));
AOI22_X1 U8751 (.B2(n11157),
.B1(REG2_REG_26__SCAN_IN),
.A1(FE_OFN8_n11821),
.A2(n12877),
.ZN(n12878));
OAI211_X1 U8752 (.C1(n13779),
.A(n12879),
.C2(n12880),
.B(n12878),
.ZN(n12881));
AOI21_X1 U8753 (.A(n12881),
.B2(FE_OFN10_n13571),
.B1(n13211),
.ZN(n12882));
OAI21_X1 U8754 (.A(n12882),
.B2(n13844),
.B1(n12883),
.ZN(n12884));
AOI21_X1 U8755 (.A(n12884),
.B2(FE_OFN9_n13503),
.B1(n12885),
.ZN(n12886));
OAI21_X1 U8756 (.A(n12886),
.B2(n13584),
.B1(n12887),
.ZN(U3264));
NAND2_X1 U8757 (.A2(n13782),
.A1(n12888),
.ZN(n12896));
AOI22_X1 U8758 (.B2(n11157),
.B1(REG2_REG_25__SCAN_IN),
.A1(FE_OFN8_n11821),
.A2(n12889),
.ZN(n12890));
OAI21_X1 U8759 (.A(n12890),
.B2(n13779),
.B1(n12891),
.ZN(n12894));
NOR2_X1 U8760 (.A2(n13844),
.A1(n12892),
.ZN(n12893));
AOI211_X1 U8761 (.C1(n13785),
.A(n12894),
.C2(n13213),
.B(n12893),
.ZN(n12895));
OAI211_X1 U8762 (.C1(n12897),
.A(n12896),
.C2(n13846),
.B(n12895),
.ZN(U3265));
NAND2_X1 U8763 (.A2(n12898),
.A1(n13029),
.ZN(n12899));
XNOR2_X1 U8764 (.B(n12899),
.A(n13030),
.ZN(n12905));
AOI21_X1 U8766 (.A(n12900),
.B2(n13655),
.B1(n13035),
.ZN(n12902));
AOI22_X1 U8767 (.B2(n13534),
.B1(n13037),
.A1(n13038),
.A2(n13689),
.ZN(n12901));
OAI211_X1 U8768 (.C1(n13041),
.A(n12902),
.C2(n12903),
.B(n12901),
.ZN(n12904));
AOI21_X1 U8769 (.A(n12904),
.B2(n13043),
.B1(n12905),
.ZN(n12906));
INV_X1 U8770 (.A(n12906),
.ZN(U3212));
INV_X1 U8771 (.A(n12942),
.ZN(n12912));
XOR2_X1 U8772 (.B(n12907),
.A(n12908),
.Z(n12911));
INV_X1 U8773 (.A(n12941),
.ZN(n12909));
NAND3_X1 U8774 (.A3(n12909),
.A1(n12912),
.A2(n12940),
.ZN(n12910));
OAI211_X1 U8775 (.C1(n12912),
.A(n12910),
.C2(n12911),
.B(n13043),
.ZN(n12916));
NOR2_X1 U8776 (.A2(STATE_REG_SCAN_IN),
.A1(n12913),
.ZN(n13319));
OAI22_X1 U8777 (.B2(n13633),
.B1(n12991),
.A1(n13427),
.A2(n13014),
.ZN(n12914));
AOI211_X1 U8778 (.C1(n13038),
.A(n13319),
.C2(n13464),
.B(n12914),
.ZN(n12915));
OAI211_X1 U8779 (.C1(n13041),
.A(n12916),
.C2(n13434),
.B(n12915),
.ZN(U3216));
AND2_X1 U8780 (.A2(n11305),
.A1(n12917),
.ZN(n12923));
INV_X1 U8781 (.A(n12918),
.ZN(n12919));
AOI21_X1 U8782 (.A(n12919),
.B2(n11305),
.B1(n12920),
.ZN(n12921));
INV_X1 U8783 (.A(n12921),
.ZN(n12922));
AOI21_X1 U8784 (.A(n12922),
.B2(n12923),
.B1(n13010),
.ZN(n12924));
INV_X1 U8785 (.A(n12924),
.ZN(n12931));
AOI22_X1 U8786 (.B2(n12932),
.B1(FE_OFN0_n11847),
.A1(n13210),
.A2(n11846),
.ZN(n12929));
AOI22_X1 U8787 (.B2(n12932),
.B1(FE_OFN22_n12925),
.A1(n13210),
.A2(FE_OFN0_n11847),
.ZN(n12927));
XNOR2_X1 U8788 (.B(FE_OFN5_n12926),
.A(n12927),
.ZN(n12928));
XOR2_X1 U8789 (.B(n12928),
.A(n12929),
.Z(n12930));
XNOR2_X1 U8790 (.B(n12930),
.A(n12931),
.ZN(n12939));
AOI22_X1 U8791 (.B2(U3149),
.B1(REG3_REG_28__SCAN_IN),
.A1(n13037),
.A2(n12932),
.ZN(n12933));
OAI21_X1 U8792 (.A(n12933),
.B2(n13041),
.B1(n12934),
.ZN(n12937));
NOR2_X1 U8793 (.A2(n12990),
.A1(n12935),
.ZN(n12936));
AOI211_X1 U8794 (.C1(n13035),
.A(n12937),
.C2(n13209),
.B(n12936),
.ZN(n12938));
OAI21_X1 U8795 (.A(n12938),
.B2(n13005),
.B1(n12939),
.ZN(U3217));
OAI21_X1 U8796 (.A(n12940),
.B2(n12941),
.B1(n12942),
.ZN(n12983));
AOI21_X1 U8797 (.A(n12984),
.B2(n12943),
.B1(n12983),
.ZN(n12947));
XNOR2_X1 U8799 (.B(n12944),
.A(n12947),
.ZN(n12953));
INV_X1 U8800 (.A(n13398),
.ZN(n12951));
OAI22_X1 U8801 (.B2(n12948),
.B1(STATE_REG_SCAN_IN),
.A1(n13427),
.A2(n12990),
.ZN(n12950));
OAI22_X1 U8802 (.B2(n13395),
.B1(n12991),
.A1(n13614),
.A2(n13014),
.ZN(n12949));
AOI211_X1 U8803 (.C1(n12951),
.A(n12950),
.C2(n13016),
.B(n12949),
.ZN(n12952));
OAI21_X1 U8804 (.A(n12952),
.B2(n13005),
.B1(n12953),
.ZN(U3220));
INV_X1 U8805 (.A(n12954),
.ZN(n12957));
INV_X1 U8806 (.A(n12955),
.ZN(n12956));
AOI21_X1 U8807 (.A(n12956),
.B2(n12957),
.B1(n13030),
.ZN(n12962));
INV_X1 U8808 (.A(n12958),
.ZN(n12960));
NAND2_X1 U8809 (.A2(n12959),
.A1(n12960),
.ZN(n12961));
XOR2_X1 U8810 (.B(n12961),
.A(n12962),
.Z(n12968));
OAI21_X1 U8811 (.A(n12963),
.B2(n13526),
.B1(n12990),
.ZN(n12964));
INV_X1 U8812 (.A(n12964),
.ZN(n12966));
AOI22_X1 U8813 (.B2(FzxTCFmmmorPYWBoKVOYVzYHHyJMkxJR_ZN),
.B1(n13037),
.A1(n13035),
.A2(n13656),
.ZN(n12965));
OAI211_X1 U8814 (.C1(n13041),
.A(n12966),
.C2(n13492),
.B(n12965),
.ZN(n12967));
AOI21_X1 U8815 (.A(n12967),
.B2(n13043),
.B1(n12968),
.ZN(n12969));
INV_X1 U8816 (.A(n12969),
.ZN(U3223));
AOI21_X1 U8817 (.A(n12970),
.B2(n12971),
.B1(n13030),
.ZN(n12975));
NAND2_X1 U8818 (.A2(n12972),
.A1(n12973),
.ZN(n12974));
XOR2_X1 U8819 (.B(n12974),
.A(n12975),
.Z(n12980));
AOI22_X1 U8820 (.B2(U3149),
.B1(REG3_REG_17__SCAN_IN),
.A1(n13035),
.A2(n13464),
.ZN(n12978));
AOI22_X1 U8821 (.B2(n12976),
.B1(n13037),
.A1(n13038),
.A2(FE_OFN6_n13667),
.ZN(n12977));
OAI211_X1 U8822 (.C1(n13041),
.A(n12978),
.C2(n13473),
.B(n12977),
.ZN(n12979));
AOI21_X1 U8823 (.A(n12979),
.B2(n13043),
.B1(n12980),
.ZN(n12981));
INV_X1 U8824 (.A(n12981),
.ZN(U3225));
XOR2_X1 U8825 (.B(n12983),
.A(n12982),
.Z(n12987));
NOR2_X1 U8826 (.A2(n12988),
.A1(n12982),
.ZN(n12985));
MUX2_X1 U8827 (.S(n12983),
.A(n12985),
.B(n12984),
.Z(n12986));
AOI21_X1 U8828 (.A(n12986),
.B2(n12987),
.B1(n12988),
.ZN(n12995));
INV_X1 U8829 (.A(n13640),
.ZN(n13456));
OAI22_X1 U8830 (.B2(n12989),
.B1(STATE_REG_SCAN_IN),
.A1(n13456),
.A2(n12990),
.ZN(n12993));
OAI22_X1 U8831 (.B2(n13407),
.B1(n12991),
.A1(n13628),
.A2(n13014),
.ZN(n12992));
AOI211_X1 U8832 (.C1(n13409),
.A(n12993),
.C2(n13016),
.B(n12992),
.ZN(n12994));
OAI21_X1 U8833 (.A(n12994),
.B2(n13005),
.B1(n12995),
.ZN(U3230));
NOR2_X1 U8834 (.A2(n12996),
.A1(n12997),
.ZN(n12999));
XOR2_X1 U8835 (.B(n12998),
.A(n12999),
.Z(n13006));
NAND2_X1 U8836 (.A2(n13214),
.A1(n13038),
.ZN(n13002));
NAND2_X1 U8837 (.A2(REG3_REG_13__SCAN_IN),
.A1(U3149),
.ZN(n13273));
NAND2_X1 U8838 (.A2(n13666),
.A1(n13035),
.ZN(n13001));
NAND2_X1 U8839 (.A2(n13554),
.A1(n13037),
.ZN(n13000));
NAND4_X1 U8840 (.A4(n13000),
.A3(n13001),
.A1(n13002),
.A2(n13273),
.ZN(n13003));
AOI21_X1 U8841 (.A(n13003),
.B2(n13551),
.B1(n13016),
.ZN(n13004));
OAI21_X1 U8842 (.A(n13004),
.B2(n13005),
.B1(n13006),
.ZN(U3231));
NAND2_X1 U8843 (.A2(n13007),
.A1(n13008),
.ZN(n13009));
XNOR2_X1 U8844 (.B(n13009),
.A(n13010),
.ZN(n13011));
NAND2_X1 U8845 (.A2(n13043),
.A1(n13011),
.ZN(n13018));
AOI22_X1 U8846 (.B2(U3149),
.B1(REG3_REG_22__SCAN_IN),
.A1(n13605),
.A2(n13038),
.ZN(n13013));
NAND2_X1 U8847 (.A2(n13604),
.A1(n13037),
.ZN(n13012));
OAI211_X1 U8848 (.C1(n13341),
.A(n13013),
.C2(n13014),
.B(n13012),
.ZN(n13015));
AOI21_X1 U8849 (.A(n13015),
.B2(n13016),
.B1(n13381),
.ZN(n13017));
NAND2_X1 U8850 (.A2(n13017),
.A1(n13018),
.ZN(U3232));
XNOR2_X1 U8851 (.B(n13019),
.A(n13020),
.ZN(n13021));
XNOR2_X1 U8852 (.B(n13021),
.A(n13022),
.ZN(n13026));
AND2_X1 U8853 (.A2(REG3_REG_18__SCAN_IN),
.A1(U3149),
.ZN(n13299));
AOI21_X1 U8854 (.A(n13299),
.B2(n13035),
.B1(n13640),
.ZN(n13024));
AOI22_X1 U8855 (.B2(n13452),
.B1(n13037),
.A1(n13038),
.A2(n13656),
.ZN(n13023));
OAI211_X1 U8856 (.C1(n13041),
.A(n13024),
.C2(n13453),
.B(n13023),
.ZN(n13025));
AOI21_X1 U8857 (.A(n13025),
.B2(n13043),
.B1(n13026),
.ZN(n13027));
INV_X1 U8858 (.A(n13027),
.ZN(U3235));
AOI21_X1 U8859 (.A(n13028),
.B2(n13029),
.B1(n13030),
.ZN(n13033));
NAND2_X1 U8860 (.A2(n13031),
.A1(n11172),
.ZN(n13032));
XOR2_X1 U8861 (.B(n13032),
.A(n13033),
.Z(n13044));
AOI21_X1 U8862 (.A(n13034),
.B2(FE_OFN6_n13667),
.B1(n13035),
.ZN(n13040));
AOI22_X1 U8863 (.B2(n13036),
.B1(n13037),
.A1(n13038),
.A2(n13666),
.ZN(n13039));
OAI211_X1 U8864 (.C1(n13041),
.A(n13040),
.C2(n13514),
.B(n13039),
.ZN(n13042));
AOI21_X1 U8865 (.A(n13042),
.B2(n13043),
.B1(n13044),
.ZN(n13045));
INV_X1 U8866 (.A(n13045),
.ZN(U3238));
INV_X1 U8870 (.A(n13208),
.ZN(n13199));
INV_X1 U8871 (.A(n13048),
.ZN(n13567));
INV_X1 U8872 (.A(n13076),
.ZN(n13050));
OAI21_X1 U8873 (.A(n13077),
.B2(n13049),
.B1(n13050),
.ZN(n13159));
AOI211_X1 U8874 (.C1(n13567),
.A(n13164),
.C2(n13157),
.B(n13159),
.ZN(n13053));
INV_X1 U8875 (.A(n13051),
.ZN(n13052));
NOR3_X1 U8876 (.A3(n13052),
.A1(n13053),
.A2(n13166),
.ZN(n13055));
NAND2_X1 U8877 (.A2(n13054),
.A1(n11227),
.ZN(n13171));
OAI21_X1 U8878 (.A(n13170),
.B2(n13171),
.B1(n13055),
.ZN(n13058));
INV_X1 U8879 (.A(n13056),
.ZN(n13057));
AOI21_X1 U8880 (.A(n13057),
.B2(n13173),
.B1(n13058),
.ZN(n13061));
NAND2_X1 U8881 (.A2(n13073),
.A1(n11182),
.ZN(n13179));
OAI21_X1 U8882 (.A(n13180),
.B2(n13179),
.B1(n13061),
.ZN(n13067));
NAND2_X1 U8883 (.A2(n13065),
.A1(n13062),
.ZN(n13063));
NOR2_X1 U8884 (.A2(n13063),
.A1(n13064),
.ZN(n13120));
OAI21_X1 U8886 (.A(n13181),
.B2(n13182),
.B1(n13066),
.ZN(n13119));
AOI21_X1 U8887 (.A(n13119),
.B2(n13120),
.B1(n13067),
.ZN(n13068));
INV_X1 U8888 (.A(n13069),
.ZN(n13198));
NOR3_X1 U8889 (.A3(n13193),
.A1(n13194),
.A2(n13198),
.ZN(n13070));
AOI21_X1 U8890 (.A(n13070),
.B2(qQydNHNCopcDTmEyGIIdyrFQIErIFgJX_ZN),
.B1(n13189),
.ZN(n13201));
INV_X1 U8891 (.A(n13071),
.ZN(n13112));
NAND2_X1 U8892 (.A2(n13072),
.A1(n13073),
.ZN(n13334));
INV_X1 U8893 (.A(n13169),
.ZN(n13349));
NOR2_X1 U8894 (.A2(n13349),
.A1(n13350),
.ZN(n13390));
INV_X1 U8895 (.A(n13170),
.ZN(n13075));
OR2_X1 U8896 (.A2(n13074),
.A1(n13075),
.ZN(n13417));
NAND2_X1 U8897 (.A2(n13076),
.A1(n13077),
.ZN(n13505));
NOR2_X1 U8898 (.A2(n13505),
.A1(n13524),
.ZN(n13079));
NAND4_X1 U8899 (.A4(n13139),
.A3(n13078),
.A1(n13421),
.A2(n13079),
.ZN(n13080));
NOR2_X1 U8900 (.A2(n13080),
.A1(n13417),
.ZN(n13081));
NAND2_X1 U8901 (.A2(n13081),
.A1(n13390),
.ZN(n13082));
NOR2_X1 U8902 (.A2(n13376),
.A1(n13082),
.ZN(n13110));
NOR2_X1 U8903 (.A2(n13083),
.A1(n13084),
.ZN(n13109));
NAND2_X1 U8905 (.A2(n13424),
.A1(n13085),
.ZN(n13467));
NAND2_X1 U8906 (.A2(n13086),
.A1(n13087),
.ZN(n13144));
NOR4_X1 U8907 (.A4(n13088),
.A3(n13144),
.A1(n13467),
.A2(n13162),
.ZN(n13107));
INV_X1 U8908 (.A(n13089),
.ZN(n13106));
NAND3_X1 U8910 (.A3(n13143),
.A1(n13092),
.A2(n13091),
.ZN(n13093));
NOR2_X1 U8911 (.A2(n13093),
.A1(n13445),
.ZN(n13105));
INV_X1 U8912 (.A(n13094),
.ZN(n13096));
AND4_X1 U8913 (.A4(n13095),
.A3(n13096),
.A1(n13098),
.A2(n13097),
.ZN(n13102));
INV_X1 U8914 (.A(n12420),
.ZN(n13101));
NOR2_X1 U8915 (.A2(n13099),
.A1(n13566),
.ZN(n13100));
AND4_X1 U8916 (.A4(n13100),
.A3(n13101),
.A1(n13920),
.A2(n13102),
.ZN(n13104));
AND4_X1 U8917 (.A4(n13104),
.A3(n13105),
.A1(n13107),
.A2(n13106),
.ZN(n13108));
NAND4_X1 U8918 (.A4(n13108),
.A3(n13109),
.A1(n13110),
.A2(n13366),
.ZN(n13111));
NOR4_X1 U8919 (.A4(n13111),
.A3(n13334),
.A1(n13113),
.A2(n13112),
.ZN(n13118));
INV_X1 U8920 (.A(n13115),
.ZN(n13116));
NAND4_X1 U8921 (.A4(n13116),
.A3(n13117),
.A1(n13118),
.A2(n12005),
.ZN(n13191));
INV_X1 U8922 (.A(n13119),
.ZN(n13188));
INV_X1 U8923 (.A(n13120),
.ZN(n13187));
INV_X1 U8924 (.A(n13121),
.ZN(n13178));
INV_X1 U8925 (.A(n13122),
.ZN(n13125));
OAI211_X1 U8926 (.C1(n13125),
.A(n13124),
.C2(n13768),
.B(n13123),
.ZN(n13127));
OAI211_X1 U8927 (.C1(FE_OFN20_n11698),
.A(n13127),
.C2(n13128),
.B(n13073),
.ZN(n13130));
OAI211_X1 U8928 (.C1(n13132),
.A(n13130),
.C2(n13131),
.B(n13129),
.ZN(n13134));
OAI211_X1 U8929 (.C1(n13221),
.A(n13134),
.C2(n13135),
.B(n13133),
.ZN(n13137));
OAI211_X1 U8930 (.C1(n13138),
.A(n13137),
.C2(n13818),
.B(n13136),
.ZN(n13142));
AOI21_X1 U8932 (.A(n13899),
.B2(n13141),
.B1(n13142),
.ZN(n13145));
OAI21_X1 U8933 (.A(n13143),
.B2(n13144),
.B1(n13145),
.ZN(n13149));
INV_X1 U8934 (.A(n13146),
.ZN(n13147));
AOI21_X1 U8935 (.A(n13147),
.B2(n13148),
.B1(n13149),
.ZN(n13152));
OAI211_X1 U8936 (.C1(n13152),
.A(n13151),
.C2(n11216),
.B(n11173),
.ZN(n13155));
NAND3_X1 U8937 (.A3(n13153),
.A1(n13155),
.A2(n13154),
.ZN(n13158));
NAND3_X1 U8938 (.A3(n13156),
.A1(n13158),
.A2(n13157),
.ZN(n13161));
INV_X1 U8939 (.A(n13159),
.ZN(n13160));
AOI21_X1 U8940 (.A(n13483),
.B2(n13160),
.B1(n13161),
.ZN(n13165));
INV_X1 U8941 (.A(n13162),
.ZN(n13163));
OAI21_X1 U8942 (.A(n13163),
.B2(n13164),
.B1(n13165),
.ZN(n13168));
AOI21_X1 U8943 (.A(n13166),
.B2(n13167),
.B1(n13168),
.ZN(n13172));
OAI211_X1 U8944 (.C1(n13172),
.A(n13170),
.C2(n13171),
.B(n13169),
.ZN(n13174));
NAND2_X1 U8945 (.A2(n13173),
.A1(n13174),
.ZN(n13176));
OAI211_X1 U8946 (.C1(n13178),
.A(n13176),
.C2(n13177),
.B(n13175),
.ZN(n13185));
NAND2_X1 U8948 (.A2(n13181),
.A1(n13182),
.ZN(n13183));
AOI21_X1 U8949 (.A(n13186),
.B2(n13187),
.B1(n13188),
.ZN(n13190));
MUX2_X1 U8950 (.S(n13189),
.A(n13191),
.B(n13190),
.Z(n13192));
OAI21_X1 U8951 (.A(n13192),
.B2(n13193),
.B1(n13194),
.ZN(n13195));
OAI21_X1 U8952 (.A(n13195),
.B2(n13196),
.B1(n13197),
.ZN(n13200));
XNOR2_X1 U8953 (.B(n13769),
.A(n13202),
.ZN(n13207));
NAND4_X1 U8954 (.A4(n13203),
.A3(n13875),
.A1(n13688),
.A2(n13204),
.ZN(n13205));
OAI211_X1 U8955 (.C1(n13767),
.A(n13205),
.C2(n13815),
.B(B_REG_SCAN_IN),
.ZN(n13206));
OAI21_X1 U8956 (.A(n13206),
.B2(n13815),
.B1(n13207),
.ZN(U3239));
MUX2_X1 U8957 (.S(n13223),
.A(n13208),
.B(DATAO_REG_31__SCAN_IN),
.Z(U3581));
MUX2_X1 U8958 (.S(U4043),
.A(DATAO_REG_29__SCAN_IN),
.B(n13209),
.Z(U3579));
MUX2_X1 U8959 (.S(U4043),
.A(DATAO_REG_28__SCAN_IN),
.B(n13210),
.Z(U3578));
MUX2_X1 U8960 (.S(U4043),
.A(DATAO_REG_27__SCAN_IN),
.B(n13211),
.Z(U3577));
MUX2_X1 U8961 (.S(U4043),
.A(DATAO_REG_26__SCAN_IN),
.B(n13212),
.Z(U3576));
MUX2_X1 U8962 (.S(U4043),
.A(DATAO_REG_25__SCAN_IN),
.B(n13343),
.Z(U3575));
MUX2_X1 U8963 (.S(U4043),
.A(DATAO_REG_24__SCAN_IN),
.B(n13213),
.Z(U3574));
MUX2_X1 U8964 (.S(U4043),
.A(DATAO_REG_23__SCAN_IN),
.B(n13587),
.Z(U3573));
MUX2_X1 U8965 (.S(U4043),
.A(DATAO_REG_22__SCAN_IN),
.B(n13362),
.Z(U3572));
MUX2_X1 U8966 (.S(U4043),
.A(DATAO_REG_21__SCAN_IN),
.B(n13605),
.Z(U3571));
MUX2_X1 U8967 (.S(U4043),
.A(DATAO_REG_20__SCAN_IN),
.B(n13612),
.Z(U3570));
MUX2_X1 U8968 (.S(U4043),
.A(DATAO_REG_19__SCAN_IN),
.B(n13640),
.Z(U3569));
MUX2_X1 U8969 (.S(U4043),
.A(DATAO_REG_18__SCAN_IN),
.B(n13464),
.Z(U3568));
MUX2_X1 U8970 (.S(U4043),
.A(DATAO_REG_17__SCAN_IN),
.B(n13656),
.Z(U3567));
MUX2_X1 U8971 (.S(U4043),
.A(DATAO_REG_16__SCAN_IN),
.B(FE_OFN6_n13667),
.Z(U3566));
MUX2_X1 U8972 (.S(U4043),
.A(DATAO_REG_15__SCAN_IN),
.B(n13655),
.Z(U3565));
MUX2_X1 U8973 (.S(U4043),
.A(DATAO_REG_14__SCAN_IN),
.B(n13666),
.Z(U3564));
MUX2_X1 U8974 (.S(U4043),
.A(DATAO_REG_13__SCAN_IN),
.B(n13689),
.Z(U3563));
MUX2_X1 U8975 (.S(U4043),
.A(DATAO_REG_12__SCAN_IN),
.B(n13214),
.Z(U3562));
MUX2_X1 U8976 (.S(U4043),
.A(DATAO_REG_11__SCAN_IN),
.B(n13687),
.Z(U3561));
MUX2_X1 U8977 (.S(U4043),
.A(DATAO_REG_10__SCAN_IN),
.B(n13215),
.Z(U3560));
MUX2_X1 U8978 (.S(n13223),
.A(n13216),
.B(DATAO_REG_9__SCAN_IN),
.Z(U3559));
MUX2_X1 U8979 (.S(U4043),
.A(DATAO_REG_8__SCAN_IN),
.B(n13217),
.Z(U3558));
MUX2_X1 U8980 (.S(U4043),
.A(DATAO_REG_7__SCAN_IN),
.B(n13218),
.Z(U3557));
MUX2_X1 U8981 (.S(U4043),
.A(DATAO_REG_6__SCAN_IN),
.B(n13219),
.Z(U3556));
MUX2_X1 U8982 (.S(U4043),
.A(DATAO_REG_5__SCAN_IN),
.B(n13220),
.Z(U3555));
MUX2_X1 U8983 (.S(n13223),
.A(n13221),
.B(DATAO_REG_4__SCAN_IN),
.Z(U3554));
MUX2_X1 U8984 (.S(U4043),
.A(DATAO_REG_3__SCAN_IN),
.B(n13784),
.Z(U3553));
MUX2_X1 U8985 (.S(n13223),
.A(FE_OFN20_n11698),
.B(DATAO_REG_2__SCAN_IN),
.Z(U3552));
MUX2_X1 U8986 (.S(U4043),
.A(DATAO_REG_1__SCAN_IN),
.B(n11358),
.Z(U3551));
MUX2_X1 U8987 (.S(n13223),
.A(n11831),
.B(DATAO_REG_0__SCAN_IN),
.Z(U3550));
AOI22_X1 U8988 (.B2(U3149),
.B1(REG3_REG_2__SCAN_IN),
.A1(FE_OFN1_n13320),
.A2(ADDR_REG_2__SCAN_IN),
.ZN(n13237));
NAND2_X1 U8989 (.A2(n13225),
.A1(n13226),
.ZN(n13231));
INV_X1 U8990 (.A(n13231),
.ZN(n13230));
NAND2_X1 U8991 (.A2(n13227),
.A1(n13228),
.ZN(n13232));
NAND2_X1 U8992 (.A2(n13232),
.A1(n13798),
.ZN(n13229));
OAI211_X1 U8993 (.C1(n13230),
.A(n13229),
.C2(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.B(n13801),
.ZN(n13234));
OAI22_X1 U8994 (.B2(n13231),
.B1(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.A1(n13795),
.A2(n13232),
.ZN(n13233));
MUX2_X1 U8995 (.S(n13777),
.A(n13234),
.B(n13233),
.Z(n13235));
INV_X1 U8996 (.A(n13235),
.ZN(n13236));
NAND3_X1 U8997 (.A3(n13236),
.A1(n13238),
.A2(n13237),
.ZN(U3242));
XNOR2_X1 U8998 (.B(REG1_REG_10__SCAN_IN),
.A(n13239),
.ZN(n13244));
INV_X1 U8999 (.A(n13244),
.ZN(n13241));
XNOR2_X1 U9000 (.B(REG2_REG_10__SCAN_IN),
.A(n13240),
.ZN(n13242));
AOI22_X1 U9001 (.B2(n13242),
.B1(n13798),
.A1(n13241),
.A2(n13804),
.ZN(n13246));
OAI21_X1 U9002 (.A(n13801),
.B2(n13242),
.B1(n13795),
.ZN(n13243));
AOI21_X1 U9003 (.A(n13243),
.B2(n13244),
.B1(n13804),
.ZN(n13245));
MUX2_X1 U9004 (.S(n13772),
.A(n13246),
.B(n13245),
.Z(n13249));
NAND2_X1 U9005 (.A2(ADDR_REG_10__SCAN_IN),
.A1(FE_OFN1_n13320),
.ZN(n13247));
NAND3_X1 U9006 (.A3(n13247),
.A1(n13249),
.A2(n13248),
.ZN(U3250));
XNOR2_X1 U9007 (.B(REG1_REG_12__SCAN_IN),
.A(n13250),
.ZN(n13252));
AOI21_X1 U9008 (.A(n13795),
.B2(n13254),
.B1(n13253),
.ZN(n13251));
AOI211_X1 U9009 (.C1(n13252),
.A(n13292),
.C2(n13804),
.B(n13251),
.ZN(n13259));
INV_X1 U9010 (.A(n13252),
.ZN(n13256));
AND2_X1 U9011 (.A2(n13798),
.A1(n13253),
.ZN(n13255));
AOI22_X1 U9012 (.B2(n13254),
.B1(n13255),
.A1(n13256),
.A2(n13804),
.ZN(n13258));
MUX2_X1 U9013 (.S(n13257),
.A(n13259),
.B(n13258),
.Z(n13262));
NAND2_X1 U9014 (.A2(ADDR_REG_12__SCAN_IN),
.A1(FE_OFN1_n13320),
.ZN(n13260));
NAND3_X1 U9015 (.A3(n13260),
.A1(n13262),
.A2(n13261),
.ZN(U3252));
XNOR2_X1 U9016 (.B(n13684),
.A(n13263),
.ZN(n13268));
INV_X1 U9017 (.A(n13268),
.ZN(n13266));
XNOR2_X1 U9018 (.B(REG2_REG_13__SCAN_IN),
.A(n13264),
.ZN(n13267));
OAI21_X1 U9019 (.A(n13801),
.B2(n13795),
.B1(n13267),
.ZN(n13265));
AOI21_X1 U9020 (.A(n13265),
.B2(n13804),
.B1(n13266),
.ZN(n13271));
AOI22_X1 U9021 (.B2(n13267),
.B1(n13798),
.A1(n13268),
.A2(n13804),
.ZN(n13270));
MUX2_X1 U9022 (.S(n13269),
.A(n13271),
.B(n13270),
.Z(n13274));
NAND2_X1 U9023 (.A2(ADDR_REG_13__SCAN_IN),
.A1(FE_OFN1_n13320),
.ZN(n13272));
NAND3_X1 U9024 (.A3(n13272),
.A1(n13274),
.A2(n13273),
.ZN(U3253));
INV_X1 U9025 (.A(n13810),
.ZN(n13812));
NOR2_X1 U9026 (.A2(n13275),
.A1(n13288),
.ZN(n13280));
NAND2_X1 U9028 (.A2(n13275),
.A1(n13288),
.ZN(n13278));
AOI21_X1 U9033 (.A(n13799),
.B2(n13794),
.B1(n13812),
.ZN(n13283));
NOR2_X1 U9034 (.A2(n13283),
.A1(REG2_REG_18__SCAN_IN),
.ZN(n13308));
INV_X1 U9035 (.A(n13308),
.ZN(n13284));
NAND2_X1 U9036 (.A2(n13283),
.A1(REG2_REG_18__SCAN_IN),
.ZN(n13306));
NAND2_X1 U9037 (.A2(NreNGPwwSfGxuZEJRmMXTmzYADEemtnb_ZN),
.A1(n13284),
.ZN(n13294));
INV_X1 U9038 (.A(n13288),
.ZN(n13285));
NAND2_X1 U9039 (.A2(REG1_REG_16__SCAN_IN),
.A1(n13285),
.ZN(n13286));
NAND2_X1 U9040 (.A2(n13663),
.A1(n13288),
.ZN(n13289));
NOR2_X1 U9041 (.A2(REG1_REG_17__SCAN_IN),
.A1(n13810),
.ZN(n13291));
XNOR2_X1 U9043 (.B(n13879),
.A(n13302),
.ZN(n13296));
NOR2_X1 U9044 (.A2(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.A1(n13296),
.ZN(n13293));
AOI211_X1 U9045 (.C1(n13294),
.A(n13293),
.C2(n13798),
.B(n13292),
.ZN(n13298));
INV_X1 U9046 (.A(n13294),
.ZN(n13295));
AOI22_X1 U9047 (.B2(n13295),
.B1(n13798),
.A1(n13296),
.A2(n13804),
.ZN(n13297));
MUX2_X1 U9048 (.S(n13307),
.A(n13298),
.B(n13297),
.Z(n13301));
AOI21_X1 U9049 (.A(n13299),
.B2(ADDR_REG_18__SCAN_IN),
.B1(FE_OFN1_n13320),
.ZN(n13300));
NAND2_X1 U9050 (.A2(n13300),
.A1(n13301),
.ZN(U3258));
XNOR2_X1 U9052 (.B(n13638),
.A(n13305),
.ZN(n13311));
OAI21_X1 U9053 (.A(NreNGPwwSfGxuZEJRmMXTmzYADEemtnb_ZN),
.B2(n13307),
.B1(n13308),
.ZN(n13309));
XNOR2_X1 U9054 (.B(REG2_REG_19__SCAN_IN),
.A(n13309),
.ZN(n13314));
OAI211_X1 U9056 (.C1(n13311),
.A(n13314),
.C2(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.B(n13801),
.ZN(n13317));
INV_X1 U9057 (.A(n13311),
.ZN(n13312));
OAI22_X1 U9058 (.B2(n13312),
.B1(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.A1(n13314),
.A2(n13795),
.ZN(n13316));
MUX2_X1 U9059 (.S(n13315),
.A(n13317),
.B(n13316),
.Z(n13318));
AOI211_X1 U9060 (.C1(FE_OFN1_n13320),
.A(n13319),
.C2(ADDR_REG_19__SCAN_IN),
.B(n13318),
.ZN(n13321));
INV_X1 U9061 (.A(n13321),
.ZN(U3259));
NAND2_X1 U9062 (.A2(n13789),
.A1(n13322),
.ZN(n13330));
INV_X1 U9063 (.A(REG2_REG_27__SCAN_IN),
.ZN(n13323));
OAI22_X1 U9064 (.B2(n13782),
.B1(n13323),
.A1(n13518),
.A2(n13324),
.ZN(n13327));
NOR2_X1 U9065 (.A2(n13844),
.A1(n13325),
.ZN(n13326));
OAI211_X1 U9066 (.C1(n13331),
.A(n13330),
.C2(n11157),
.B(n13329),
.ZN(U3263));
XOR2_X1 U9067 (.B(n13332),
.A(n13334),
.Z(n13592));
INV_X1 U9068 (.A(n13592),
.ZN(n13347));
XNOR2_X1 U9069 (.B(n13334),
.A(n13333),
.ZN(n13585));
INV_X1 U9071 (.A(n12139),
.ZN(n13336));
OAI21_X1 U9072 (.A(n13336),
.B2(n13337),
.B1(n11798),
.ZN(n13709));
AOI22_X1 U9073 (.B2(n11157),
.B1(REG2_REG_24__SCAN_IN),
.A1(FE_OFN8_n11821),
.A2(n13586),
.ZN(n13340));
NAND2_X1 U9074 (.A2(n13842),
.A1(n13338),
.ZN(n13339));
OAI211_X1 U9075 (.C1(n13341),
.A(n13340),
.C2(n13577),
.B(n13339),
.ZN(n13342));
AOI21_X1 U9076 (.A(n13342),
.B2(FE_OFN10_n13571),
.B1(n13343),
.ZN(n13344));
OAI21_X1 U9077 (.A(n13344),
.B2(n13844),
.B1(n13709),
.ZN(n13345));
AOI21_X1 U9078 (.A(n13345),
.B2(n13585),
.B1(FE_OFN9_n13503),
.ZN(n13346));
OAI21_X1 U9079 (.A(n13346),
.B2(n13584),
.B1(n13347),
.ZN(U3266));
NAND2_X1 U9084 (.A2(n13353),
.A1(n13379),
.ZN(n13354));
XNOR2_X1 U9085 (.B(n13366),
.A(n13354),
.ZN(n13357));
NOR2_X1 U9086 (.A2(n13627),
.A1(n13355),
.ZN(n13356));
AOI21_X1 U9087 (.A(n11798),
.B2(n13358),
.B1(n13360),
.ZN(n13712));
AOI22_X1 U9088 (.B2(n11157),
.B1(REG2_REG_23__SCAN_IN),
.A1(n13361),
.A2(n13842),
.ZN(n13364));
NAND2_X1 U9089 (.A2(n13785),
.A1(n13362),
.ZN(n13363));
OAI211_X1 U9090 (.C1(n13518),
.A(n13364),
.C2(n13595),
.B(n13363),
.ZN(n13370));
NOR2_X1 U9093 (.A2(n13584),
.A1(n13598),
.ZN(n13369));
AOI211_X1 U9094 (.C1(n13712),
.A(n13370),
.C2(FE_OFN2_n13580),
.B(n13369),
.ZN(n13371));
OAI21_X1 U9095 (.A(n13371),
.B2(n13601),
.B1(n11157),
.ZN(U3267));
XNOR2_X1 U9096 (.B(n13376),
.A(n13372),
.ZN(n13606));
INV_X1 U9097 (.A(n13606),
.ZN(n13388));
OAI211_X1 U9098 (.C1(n13373),
.A(n13358),
.C2(n13384),
.B(n13374),
.ZN(n13607));
NAND3_X1 U9099 (.A3(n13375),
.A1(n13377),
.A2(n13376),
.ZN(n13378));
AOI21_X1 U9100 (.A(n13568),
.B2(n13378),
.B1(n13379),
.ZN(n13380));
AOI21_X1 U9101 (.A(n13380),
.B2(n13587),
.B1(n13690),
.ZN(n13610));
OAI21_X1 U9102 (.A(n13610),
.B2(n13607),
.B1(n13769),
.ZN(n13386));
AOI22_X1 U9103 (.B2(n11157),
.B1(REG2_REG_22__SCAN_IN),
.A1(n13381),
.A2(n13842),
.ZN(n13383));
NAND2_X1 U9104 (.A2(n13785),
.A1(n13605),
.ZN(n13382));
OAI211_X1 U9105 (.C1(n13518),
.A(n13383),
.C2(n13384),
.B(n13382),
.ZN(n13385));
AOI21_X1 U9106 (.A(n13385),
.B2(n13782),
.B1(n13386),
.ZN(n13387));
OAI21_X1 U9107 (.A(n13387),
.B2(n13388),
.B1(n13584),
.ZN(U3268));
INV_X1 U9108 (.A(n13390),
.ZN(n13391));
XNOR2_X1 U9109 (.B(n13391),
.A(n13389),
.ZN(n13620));
XNOR2_X1 U9110 (.B(n13391),
.A(n13348),
.ZN(n13616));
NOR2_X1 U9111 (.A2(n13395),
.A1(n13392),
.ZN(n13393));
OR2_X1 U9112 (.A2(n13393),
.A1(n13373),
.ZN(n13718));
INV_X1 U9113 (.A(FE_OFN10_n13571),
.ZN(n13455));
OAI22_X1 U9114 (.B2(n13395),
.B1(n13518),
.A1(n13614),
.A2(n13455),
.ZN(n13400));
NAND2_X1 U9115 (.A2(n13785),
.A1(n13612),
.ZN(n13397));
NAND2_X1 U9116 (.A2(REG2_REG_21__SCAN_IN),
.A1(n11157),
.ZN(n13396));
OAI211_X1 U9117 (.C1(n13779),
.A(n13397),
.C2(n13398),
.B(rlUqTqnDczmjZLOdxrCVPPbsubqicwLv_Z),
.ZN(n13399));
NOR2_X1 U9118 (.A2(n13399),
.A1(n13400),
.ZN(n13401));
OAI21_X1 U9119 (.A(n13401),
.B2(n13844),
.B1(n13718),
.ZN(n13402));
OR3_X1 U9120 (.A3(n13616),
.A2(n13402),
.A1(FE_OFN9_n13503),
.ZN(n13403));
OAI21_X1 U9121 (.A(n13403),
.B2(n13620),
.B1(n13584),
.ZN(U3269));
NOR2_X1 U9124 (.A2(n13407),
.A1(n13406),
.ZN(n13408));
OR2_X1 U9125 (.A2(n13408),
.A1(n13392),
.ZN(n13722));
INV_X1 U9126 (.A(n13722),
.ZN(n13415));
NAND2_X1 U9127 (.A2(FE_OFN10_n13571),
.A1(n13605),
.ZN(n13413));
AOI22_X1 U9128 (.B2(REG2_REG_20__SCAN_IN),
.B1(n11157),
.A1(n13409),
.A2(n13842),
.ZN(n13412));
NAND2_X1 U9129 (.A2(n13640),
.A1(n13785),
.ZN(n13411));
NAND2_X1 U9130 (.A2(n13624),
.A1(FE_OFN8_n11821),
.ZN(n13410));
NAND4_X1 U9131 (.A4(n13410),
.A3(n13411),
.A1(n13413),
.A2(n13412),
.ZN(n13414));
AOI21_X1 U9132 (.A(n13414),
.B2(FE_OFN2_n13580),
.B1(n13415),
.ZN(n13419));
XNOR2_X1 U9133 (.B(n13417),
.A(n13416),
.ZN(n13630));
NAND2_X1 U9134 (.A2(n13789),
.A1(n13630),
.ZN(n13418));
OAI211_X1 U9135 (.C1(n13626),
.A(n13419),
.C2(n11157),
.B(n13418),
.ZN(U3270));
OAI21_X1 U9139 (.A(n13443),
.B2(n13445),
.B1(n13446),
.ZN(n13426));
XOR2_X1 U9140 (.B(n13426),
.A(n13430),
.Z(n13428));
OAI22_X1 U9141 (.B2(n13627),
.B1(n13427),
.A1(n13428),
.A2(n13568),
.ZN(n13635));
INV_X1 U9142 (.A(n13635),
.ZN(n13442));
INV_X1 U9144 (.A(n13406),
.ZN(n13433));
NAND2_X1 U9147 (.A2(n13432),
.A1(n13433),
.ZN(n13726));
INV_X1 U9148 (.A(n13464),
.ZN(n13634));
INV_X1 U9149 (.A(n13434),
.ZN(n13435));
AOI22_X1 U9150 (.B2(n13435),
.B1(n13842),
.A1(n11157),
.A2(REG2_REG_19__SCAN_IN),
.ZN(n13436));
OAI21_X1 U9151 (.A(n13436),
.B2(n13634),
.B1(n13577),
.ZN(n13437));
AOI21_X1 U9152 (.A(n13437),
.B2(FE_OFN8_n11821),
.B1(n13438),
.ZN(n13439));
OAI21_X1 U9153 (.A(n13439),
.B2(n13844),
.B1(n13726),
.ZN(n13440));
AOI21_X1 U9154 (.A(n13440),
.B2(n13789),
.B1(n13637),
.ZN(n13441));
OAI21_X1 U9155 (.A(n13441),
.B2(n11157),
.B1(n13442),
.ZN(U3271));
INV_X1 U9156 (.A(n13443),
.ZN(n13444));
NOR2_X1 U9157 (.A2(n13444),
.A1(n13445),
.ZN(n13448));
XNOR2_X1 U9158 (.B(n13448),
.A(n13446),
.ZN(n13447));
NAND2_X1 U9159 (.A2(n13672),
.A1(n13447),
.ZN(n13647));
NAND3_X1 U9162 (.A3(n13431),
.A1(n13452),
.A2(n13470),
.ZN(n13730));
INV_X1 U9163 (.A(n13730),
.ZN(n13460));
OAI22_X1 U9164 (.B2(n13779),
.B1(n13453),
.A1(n13782),
.A2(n13454),
.ZN(n13458));
OAI22_X1 U9165 (.B2(n13643),
.B1(n13518),
.A1(n13456),
.A2(n13455),
.ZN(n13457));
AOI211_X1 U9166 (.C1(n13785),
.A(n13458),
.C2(n13656),
.B(n13457),
.ZN(n13459));
OAI21_X1 U9167 (.A(n13459),
.B2(n13844),
.B1(n13460),
.ZN(n13461));
AOI21_X1 U9168 (.A(n13461),
.B2(n13645),
.B1(n13789),
.ZN(n13462));
OAI21_X1 U9169 (.A(n13462),
.B2(n11157),
.B1(n13647),
.ZN(U3272));
XNOR2_X1 U9170 (.B(n13467),
.A(n13422),
.ZN(n13463));
NAND2_X1 U9171 (.A2(n13672),
.A1(n13463),
.ZN(n13466));
AOI22_X1 U9172 (.B2(FE_OFN6_n13667),
.B1(n13688),
.A1(n13464),
.A2(n13690),
.ZN(n13465));
OAI211_X1 U9173 (.C1(n13698),
.A(n13466),
.C2(n13471),
.B(n13465),
.ZN(n13651));
INV_X1 U9174 (.A(n13651),
.ZN(n13478));
XNOR2_X1 U9175 (.B(n13467),
.A(n13468),
.ZN(n13652));
INV_X1 U9176 (.A(n13469),
.ZN(n13472));
OAI21_X1 U9177 (.A(n13470),
.B2(n13471),
.B1(n13472),
.ZN(n13735));
INV_X1 U9178 (.A(n13473),
.ZN(n13474));
AOI22_X1 U9179 (.B2(n13474),
.B1(n13842),
.A1(n11157),
.A2(REG2_REG_17__SCAN_IN),
.ZN(n13475));
OAI21_X1 U9180 (.A(n13475),
.B2(n13844),
.B1(n13735),
.ZN(n13476));
AOI21_X1 U9181 (.A(n13476),
.B2(n13789),
.B1(n13652),
.ZN(n13477));
OAI21_X1 U9182 (.A(n13477),
.B2(n11157),
.B1(n13478),
.ZN(U3273));
OAI21_X1 U9183 (.A(n13479),
.B2(n13486),
.B1(n13480),
.ZN(n13661));
INV_X1 U9184 (.A(n13661),
.ZN(n13500));
OAI21_X1 U9185 (.A(n13482),
.B2(n13483),
.B1(n11234),
.ZN(n13502));
INV_X1 U9186 (.A(n13484),
.ZN(n13509));
NAND2_X1 U9187 (.A2(n13509),
.A1(n13502),
.ZN(n13501));
NAND2_X1 U9188 (.A2(n13485),
.A1(n13501),
.ZN(n13487));
XNOR2_X1 U9189 (.B(n13486),
.A(n13487),
.ZN(n13489));
OAI22_X1 U9190 (.B2(n13488),
.B1(n13500),
.A1(n13489),
.A2(n13568),
.ZN(n13659));
NAND2_X1 U9191 (.A2(n13782),
.A1(n13659),
.ZN(n13499));
OAI21_X1 U9192 (.A(n13469),
.B2(n13658),
.B1(n13490),
.ZN(n13739));
INV_X1 U9193 (.A(n13739),
.ZN(n13497));
AOI22_X1 U9194 (.B2(n13656),
.B1(FE_OFN10_n13571),
.A1(FzxTCFmmmorPYWBoKVOYVzYHHyJMkxJR_ZN),
.A2(FE_OFN8_n11821),
.ZN(n13495));
INV_X1 U9195 (.A(n13492),
.ZN(n13493));
AOI22_X1 U9196 (.B2(n13493),
.B1(n13842),
.A1(n11157),
.A2(REG2_REG_16__SCAN_IN),
.ZN(n13494));
OAI211_X1 U9197 (.C1(n13526),
.A(n13495),
.C2(n13577),
.B(n13494),
.ZN(n13496));
AOI21_X1 U9198 (.A(n13496),
.B2(FE_OFN2_n13580),
.B1(n13497),
.ZN(n13498));
OAI211_X1 U9199 (.C1(n13500),
.A(n13499),
.C2(n13846),
.B(n13498),
.ZN(U3274));
OAI21_X1 U9200 (.A(n13501),
.B2(n13509),
.B1(n13502),
.ZN(n13673));
INV_X1 U9201 (.A(n13673),
.ZN(n13523));
INV_X1 U9202 (.A(FE_OFN9_n13503),
.ZN(n13522));
NAND2_X1 U9203 (.A2(n13506),
.A1(n13507),
.ZN(n13531));
INV_X1 U9204 (.A(n13524),
.ZN(n13530));
INV_X1 U9206 (.A(n13508),
.ZN(n13510));
OAI21_X1 U9207 (.A(n13509),
.B2(n13510),
.B1(n13533),
.ZN(n13512));
NAND2_X1 U9208 (.A2(n13511),
.A1(n13512),
.ZN(n13665));
INV_X1 U9209 (.A(n13490),
.ZN(n13513));
OAI21_X1 U9210 (.A(n13513),
.B2(n13670),
.B1(n13535),
.ZN(n13743));
NOR2_X1 U9211 (.A2(n13844),
.A1(n13743),
.ZN(n13520));
AOI22_X1 U9212 (.B2(FE_OFN6_n13667),
.B1(FE_OFN10_n13571),
.A1(n13785),
.A2(n13666),
.ZN(n13517));
INV_X1 U9213 (.A(n13514),
.ZN(n13515));
AOI22_X1 U9214 (.B2(n13515),
.B1(n13842),
.A1(n11157),
.A2(REG2_REG_15__SCAN_IN),
.ZN(n13516));
OAI211_X1 U9215 (.C1(n13670),
.A(n13517),
.C2(n13518),
.B(n13516),
.ZN(n13519));
AOI211_X1 U9216 (.C1(n13665),
.A(n13520),
.C2(n13789),
.B(n13519),
.ZN(n13521));
OAI21_X1 U9217 (.A(n13521),
.B2(n13522),
.B1(n13523),
.ZN(U3275));
XNOR2_X1 U9218 (.B(n13524),
.A(n13481),
.ZN(n13529));
OAI22_X1 U9219 (.B2(n13525),
.B1(n13819),
.A1(n13526),
.A2(n13627),
.ZN(n13527));
AOI21_X1 U9220 (.A(n13527),
.B2(n13623),
.B1(n13534),
.ZN(n13528));
OAI21_X1 U9221 (.A(n13528),
.B2(n13568),
.B1(n13529),
.ZN(n13675));
INV_X1 U9222 (.A(n13675),
.ZN(n13541));
AND2_X1 U9225 (.A2(n13534),
.A1(n13550),
.ZN(n13536));
OR2_X1 U9226 (.A2(n13535),
.A1(n13536),
.ZN(n13747));
AOI22_X1 U9227 (.B2(n13537),
.B1(n13842),
.A1(n11157),
.A2(REG2_REG_14__SCAN_IN),
.ZN(n13538));
OAI21_X1 U9228 (.A(n13538),
.B2(n13844),
.B1(n13747),
.ZN(n13539));
AOI21_X1 U9229 (.A(n13539),
.B2(n13789),
.B1(n13676),
.ZN(n13540));
OAI21_X1 U9230 (.A(n13540),
.B2(n11157),
.B1(n13541),
.ZN(U3276));
NAND2_X1 U9231 (.A2(n13542),
.A1(n13543),
.ZN(n13544));
XNOR2_X1 U9232 (.B(n13547),
.A(n13544),
.ZN(n13546));
OAI22_X1 U9233 (.B2(n13627),
.B1(n13545),
.A1(n13546),
.A2(n13568),
.ZN(n13681));
INV_X1 U9234 (.A(n13681),
.ZN(n13558));
XNOR2_X1 U9235 (.B(n13547),
.A(n13504),
.ZN(n13683));
NAND2_X1 U9236 (.A2(n13554),
.A1(n13548),
.ZN(n13549));
NAND2_X1 U9237 (.A2(n13549),
.A1(n13550),
.ZN(n13751));
AOI22_X1 U9238 (.B2(n13551),
.B1(n13842),
.A1(n11157),
.A2(REG2_REG_13__SCAN_IN),
.ZN(n13552));
OAI21_X1 U9239 (.A(n13552),
.B2(n13680),
.B1(n13577),
.ZN(n13553));
AOI21_X1 U9240 (.A(n13553),
.B2(FE_OFN8_n11821),
.B1(n13554),
.ZN(n13555));
OAI21_X1 U9241 (.A(n13555),
.B2(n13844),
.B1(n13751),
.ZN(n13556));
AOI21_X1 U9242 (.A(n13556),
.B2(n13789),
.B1(n13683),
.ZN(n13557));
OAI21_X1 U9243 (.A(n13557),
.B2(n11157),
.B1(n13558),
.ZN(U3277));
NAND2_X1 U9244 (.A2(n13559),
.A1(n12686),
.ZN(n13563));
AND2_X1 U9245 (.A2(n13563),
.A1(n13561),
.ZN(n13565));
NAND2_X1 U9246 (.A2(n13562),
.A1(n13563),
.ZN(n13564));
OAI21_X1 U9247 (.A(n13564),
.B2(n13566),
.B1(n13565),
.ZN(n13686));
XNOR2_X1 U9248 (.B(n13566),
.A(n13567),
.ZN(n13569));
NOR2_X1 U9249 (.A2(n13568),
.A1(n13569),
.ZN(n13693));
NAND2_X1 U9250 (.A2(n13782),
.A1(n13693),
.ZN(n13583));
OAI21_X1 U9251 (.A(n13548),
.B2(n13692),
.B1(n13570),
.ZN(n13755));
INV_X1 U9252 (.A(n13755),
.ZN(n13581));
AOI22_X1 U9253 (.B2(n13689),
.B1(FE_OFN10_n13571),
.A1(n13572),
.A2(FE_OFN8_n11821),
.ZN(n13576));
INV_X1 U9254 (.A(n13573),
.ZN(n13574));
AOI22_X1 U9255 (.B2(n13574),
.B1(n13842),
.A1(n11157),
.A2(REG2_REG_12__SCAN_IN),
.ZN(n13575));
OAI211_X1 U9256 (.C1(n13578),
.A(n13576),
.C2(n13577),
.B(n13575),
.ZN(n13579));
AOI21_X1 U9257 (.A(n13579),
.B2(FE_OFN2_n13580),
.B1(n13581),
.ZN(n13582));
OAI211_X1 U9258 (.C1(n13584),
.A(n13583),
.C2(n13686),
.B(n13582),
.ZN(U3278));
NAND2_X1 U9259 (.A2(n13672),
.A1(n13585),
.ZN(n13589));
AOI22_X1 U9260 (.B2(n13586),
.B1(n13623),
.A1(n13587),
.A2(n13688),
.ZN(n13588));
OAI211_X1 U9261 (.C1(n13890),
.A(n13589),
.C2(n13627),
.B(n13588),
.ZN(n13591));
AOI21_X1 U9262 (.A(n13591),
.B2(n13829),
.B1(n13592),
.ZN(n13706));
MUX2_X1 U9263 (.S(n13841),
.A(n13593),
.B(n13706),
.Z(n13594));
OAI21_X1 U9264 (.A(n13594),
.B2(n13709),
.B1(FE_OFN7_n13835),
.ZN(U3542));
OAI22_X1 U9265 (.B2(n13698),
.B1(n13595),
.A1(n13614),
.A2(n13819),
.ZN(n13596));
NAND2_X1 U9267 (.A2(n13600),
.A1(n13601),
.ZN(n13710));
MUX2_X1 U9268 (.S(n13841),
.A(REG1_REG_23__SCAN_IN),
.B(n13710),
.Z(n13602));
AOI21_X1 U9269 (.A(n13602),
.B2(n13712),
.B1(n13649),
.ZN(n13603));
INV_X1 U9270 (.A(n13603),
.ZN(U3541));
AOI22_X1 U9271 (.B2(n13623),
.B1(n13604),
.A1(n13605),
.A2(n13688),
.ZN(n13609));
NAND2_X1 U9272 (.A2(n13829),
.A1(n13606),
.ZN(n13608));
NAND4_X1 U9273 (.A4(n13607),
.A3(n13608),
.A1(n13610),
.A2(n13609),
.ZN(n13714));
MUX2_X1 U9274 (.S(n13841),
.A(REG1_REG_22__SCAN_IN),
.B(n13714),
.Z(U3540));
AOI22_X1 U9275 (.B2(n13623),
.B1(n13611),
.A1(n13612),
.A2(n13688),
.ZN(n13613));
OAI21_X1 U9276 (.A(n13613),
.B2(n13627),
.B1(n13614),
.ZN(n13615));
INV_X1 U9277 (.A(n13615),
.ZN(n13618));
NAND2_X1 U9278 (.A2(n13672),
.A1(n13616),
.ZN(n13617));
OAI211_X1 U9279 (.C1(n13620),
.A(n13618),
.C2(n13619),
.B(n13617),
.ZN(n13715));
MUX2_X1 U9280 (.S(n13841),
.A(REG1_REG_21__SCAN_IN),
.B(n13715),
.Z(n13621));
INV_X1 U9281 (.A(n13621),
.ZN(n13622));
OAI21_X1 U9282 (.A(n13622),
.B2(n13718),
.B1(FE_OFN7_n13835),
.ZN(U3539));
AOI22_X1 U9283 (.B2(n13623),
.B1(n13624),
.A1(n13640),
.A2(n13688),
.ZN(n13625));
OAI211_X1 U9284 (.C1(n13628),
.A(n13626),
.C2(n13627),
.B(n13625),
.ZN(n13629));
AOI21_X1 U9285 (.A(n13629),
.B2(n13630),
.B1(n13829),
.ZN(n13719));
MUX2_X1 U9286 (.S(n13841),
.A(n13631),
.B(n13719),
.Z(n13632));
OAI21_X1 U9287 (.A(n13632),
.B2(n13722),
.B1(FE_OFN7_n13835),
.ZN(U3538));
OAI22_X1 U9288 (.B2(n13698),
.B1(n13633),
.A1(n13634),
.A2(n13819),
.ZN(n13636));
AOI211_X1 U9289 (.C1(n13637),
.A(n13636),
.C2(n13829),
.B(n13635),
.ZN(n13723));
MUX2_X1 U9290 (.S(n13841),
.A(n13638),
.B(n13723),
.Z(n13639));
OAI21_X1 U9291 (.A(n13639),
.B2(n13726),
.B1(FE_OFN7_n13835),
.ZN(U3537));
NAND2_X1 U9292 (.A2(n13690),
.A1(n13640),
.ZN(n13642));
NAND2_X1 U9293 (.A2(n13688),
.A1(n13656),
.ZN(n13641));
OAI211_X1 U9294 (.C1(n13698),
.A(n13642),
.C2(n13643),
.B(n13641),
.ZN(n13644));
AOI21_X1 U9295 (.A(n13644),
.B2(n13829),
.B1(n13645),
.ZN(n13646));
NAND2_X1 U9296 (.A2(n13646),
.A1(n13647),
.ZN(n13727));
MUX2_X1 U9297 (.S(n13839),
.A(n13727),
.B(REG1_REG_18__SCAN_IN),
.Z(n13648));
AOI21_X1 U9298 (.A(n13648),
.B2(n13730),
.B1(n13649),
.ZN(n13650));
INV_X1 U9299 (.A(n13650),
.ZN(U3536));
AOI21_X1 U9300 (.A(n13651),
.B2(n13652),
.B1(n13829),
.ZN(n13732));
MUX2_X1 U9301 (.S(n13841),
.A(n13653),
.B(n13732),
.Z(n13654));
OAI21_X1 U9302 (.A(n13654),
.B2(n13735),
.B1(FE_OFN7_n13835),
.ZN(U3535));
AOI22_X1 U9303 (.B2(n13688),
.B1(n13655),
.A1(n13656),
.A2(n13690),
.ZN(n13657));
OAI21_X1 U9304 (.A(n13657),
.B2(n13698),
.B1(n13658),
.ZN(n13660));
AOI211_X1 U9305 (.C1(n13662),
.A(n13660),
.C2(n13661),
.B(n13659),
.ZN(n13736));
MUX2_X1 U9306 (.S(n13841),
.A(n13663),
.B(n13736),
.Z(n13664));
OAI21_X1 U9307 (.A(n13664),
.B2(n13739),
.B1(FE_OFN7_n13835),
.ZN(U3534));
NAND2_X1 U9308 (.A2(n13829),
.A1(n13665),
.ZN(n13669));
AOI22_X1 U9309 (.B2(n13666),
.B1(n13688),
.A1(n13690),
.A2(FE_OFN6_n13667),
.ZN(n13668));
OAI211_X1 U9310 (.C1(n13698),
.A(n13669),
.C2(n13670),
.B(n13668),
.ZN(n13671));
AOI21_X1 U9311 (.A(n13671),
.B2(n13672),
.B1(n13673),
.ZN(n13740));
MUX2_X1 U9312 (.S(n13841),
.A(n12772),
.B(n13740),
.Z(n13674));
OAI21_X1 U9313 (.A(n13674),
.B2(n13743),
.B1(FE_OFN7_n13835),
.ZN(U3533));
INV_X1 U9314 (.A(REG1_REG_14__SCAN_IN),
.ZN(n13677));
AOI21_X1 U9315 (.A(n13675),
.B2(n13829),
.B1(n13676),
.ZN(n13744));
MUX2_X1 U9316 (.S(n13841),
.A(n13677),
.B(n13744),
.Z(n13678));
OAI21_X1 U9317 (.A(n13678),
.B2(n13747),
.B1(FE_OFN7_n13835),
.ZN(U3532));
OAI22_X1 U9318 (.B2(n13679),
.B1(n13698),
.A1(n13819),
.A2(n13680),
.ZN(n13682));
AOI211_X1 U9319 (.C1(n13683),
.A(n13682),
.C2(n13829),
.B(n13681),
.ZN(n13748));
MUX2_X1 U9320 (.S(n13841),
.A(n13684),
.B(n13748),
.Z(n13685));
OAI21_X1 U9321 (.A(n13685),
.B2(n13751),
.B1(FE_OFN7_n13835),
.ZN(U3531));
INV_X1 U9322 (.A(n13686),
.ZN(n13695));
AOI22_X1 U9323 (.B2(n13687),
.B1(n13688),
.A1(n13690),
.A2(n13689),
.ZN(n13691));
OAI21_X1 U9324 (.A(n13691),
.B2(n13698),
.B1(n13692),
.ZN(n13694));
AOI211_X1 U9325 (.C1(n13695),
.A(n13694),
.C2(n13829),
.B(n13693),
.ZN(n13752));
MUX2_X1 U9326 (.S(n13841),
.A(n13696),
.B(n13752),
.Z(n13697));
OAI21_X1 U9327 (.A(n13697),
.B2(n13755),
.B1(FE_OFN7_n13835),
.ZN(U3530));
OAI22_X1 U9328 (.B2(n13698),
.B1(n13699),
.A1(n13819),
.A2(n13700),
.ZN(n13702));
AOI211_X1 U9329 (.C1(n13703),
.A(n13702),
.C2(n13829),
.B(n13701),
.ZN(n13756));
MUX2_X1 U9330 (.S(n13841),
.A(n13704),
.B(n13756),
.Z(n13705));
OAI21_X1 U9331 (.A(n13705),
.B2(n13760),
.B1(FE_OFN7_n13835),
.ZN(U3529));
INV_X1 U9332 (.A(REG0_REG_24__SCAN_IN),
.ZN(n13707));
MUX2_X1 U9333 (.S(FE_OFN3_n13832),
.A(n13707),
.B(n13706),
.Z(n13708));
OAI21_X1 U9334 (.A(n13708),
.B2(FE_OFN21_n13759),
.B1(n13709),
.ZN(U3510));
MUX2_X1 U9335 (.S(FE_OFN3_n13832),
.A(REG0_REG_23__SCAN_IN),
.B(n13710),
.Z(n13711));
AOI21_X1 U9336 (.A(n13711),
.B2(n13729),
.B1(n13712),
.ZN(n13713));
INV_X1 U9337 (.A(n13713),
.ZN(U3509));
MUX2_X1 U9338 (.S(FE_OFN3_n13832),
.A(REG0_REG_22__SCAN_IN),
.B(n13714),
.Z(U3508));
MUX2_X1 U9339 (.S(FE_OFN3_n13832),
.A(REG0_REG_21__SCAN_IN),
.B(n13715),
.Z(n13716));
INV_X1 U9340 (.A(n13716),
.ZN(n13717));
OAI21_X1 U9341 (.A(n13717),
.B2(FE_OFN21_n13759),
.B1(n13718),
.ZN(U3507));
INV_X1 U9342 (.A(REG0_REG_20__SCAN_IN),
.ZN(n13720));
MUX2_X1 U9343 (.S(FE_OFN3_n13832),
.A(n13720),
.B(n13719),
.Z(n13721));
OAI21_X1 U9344 (.A(n13721),
.B2(FE_OFN21_n13759),
.B1(n13722),
.ZN(U3506));
INV_X1 U9345 (.A(REG0_REG_19__SCAN_IN),
.ZN(n13724));
MUX2_X1 U9346 (.S(FE_OFN3_n13832),
.A(n13724),
.B(n13723),
.Z(n13725));
OAI21_X1 U9347 (.A(n13725),
.B2(FE_OFN21_n13759),
.B1(n13726),
.ZN(U3505));
MUX2_X1 U9348 (.S(n13860),
.A(n13727),
.B(REG0_REG_18__SCAN_IN),
.Z(n13728));
AOI21_X1 U9349 (.A(n13728),
.B2(n13729),
.B1(n13730),
.ZN(n13731));
INV_X1 U9350 (.A(n13731),
.ZN(U3503));
INV_X1 U9351 (.A(REG0_REG_17__SCAN_IN),
.ZN(n13733));
MUX2_X1 U9352 (.S(FE_OFN3_n13832),
.A(n13733),
.B(n13732),
.Z(n13734));
OAI21_X1 U9353 (.A(n13734),
.B2(FE_OFN21_n13759),
.B1(n13735),
.ZN(U3501));
INV_X1 U9354 (.A(REG0_REG_16__SCAN_IN),
.ZN(n12805));
MUX2_X1 U9355 (.S(FE_OFN3_n13832),
.A(n13737),
.B(n13736),
.Z(n13738));
OAI21_X1 U9356 (.A(n13738),
.B2(FE_OFN21_n13759),
.B1(n13739),
.ZN(U3499));
INV_X1 U9357 (.A(REG0_REG_15__SCAN_IN),
.ZN(n13741));
MUX2_X1 U9358 (.S(FE_OFN3_n13832),
.A(n13741),
.B(n13740),
.Z(n13742));
OAI21_X1 U9359 (.A(n13742),
.B2(FE_OFN21_n13759),
.B1(n13743),
.ZN(U3497));
MUX2_X1 U9360 (.S(FE_OFN3_n13832),
.A(n13745),
.B(n13744),
.Z(n13746));
OAI21_X1 U9361 (.A(n13746),
.B2(FE_OFN21_n13759),
.B1(n13747),
.ZN(U3495));
MUX2_X1 U9362 (.S(FE_OFN3_n13832),
.A(n13749),
.B(n13748),
.Z(n13750));
OAI21_X1 U9363 (.A(n13750),
.B2(FE_OFN21_n13759),
.B1(n13751),
.ZN(U3493));
MUX2_X1 U9364 (.S(FE_OFN3_n13832),
.A(n13753),
.B(n13752),
.Z(n13754));
OAI21_X1 U9365 (.A(n13754),
.B2(FE_OFN21_n13759),
.B1(n13755),
.ZN(U3491));
MUX2_X1 U9366 (.S(FE_OFN3_n13832),
.A(n13757),
.B(n13756),
.Z(n13758));
OAI21_X1 U9367 (.A(n13758),
.B2(FE_OFN21_n13759),
.B1(n13760),
.ZN(U3489));
MUX2_X1 U9368 (.S(n13814),
.A(n13761),
.B(D_REG_1__SCAN_IN),
.Z(U3459));
MUX2_X1 U9369 (.S(U3149),
.A(n13762),
.B(DATAI_30_),
.Z(U3322));
MUX2_X1 U9370 (.S(U3149),
.A(n13763),
.B(DATAI_29_),
.Z(U3323));
MUX2_X1 U9371 (.S(STATE_REG_SCAN_IN),
.A(DATAI_28_),
.B(n13764),
.Z(U3324));
MUX2_X1 U9372 (.S(STATE_REG_SCAN_IN),
.A(DATAI_27_),
.B(n13875),
.Z(U3325));
MUX2_X1 U9373 (.S(U3149),
.A(n13766),
.B(DATAI_26_),
.Z(U3326));
MUX2_X1 U9374 (.S(STATE_REG_SCAN_IN),
.A(DATAI_22_),
.B(n13767),
.Z(U3330));
MUX2_X1 U9375 (.S(U3149),
.A(n13768),
.B(DATAI_21_),
.Z(U3331));
MUX2_X1 U9376 (.S(STATE_REG_SCAN_IN),
.A(DATAI_20_),
.B(n11244),
.Z(U3332));
MUX2_X1 U9377 (.S(U3149),
.A(n13769),
.B(DATAI_19_),
.Z(U3333));
MUX2_X1 U9378 (.S(U3149),
.A(n13770),
.B(DATAI_14_),
.Z(U3338));
MUX2_X1 U9379 (.S(U3149),
.A(n13771),
.B(DATAI_11_),
.Z(U3341));
MUX2_X1 U9380 (.S(STATE_REG_SCAN_IN),
.A(DATAI_10_),
.B(n13772),
.Z(U3342));
MUX2_X1 U9381 (.S(U3149),
.A(n13773),
.B(DATAI_9_),
.Z(U3343));
MUX2_X1 U9382 (.S(U3149),
.A(n13774),
.B(DATAI_6_),
.Z(U3346));
MUX2_X1 U9383 (.S(U3149),
.A(n13775),
.B(DATAI_5_),
.Z(U3347));
MUX2_X1 U9384 (.S(U3149),
.A(n13776),
.B(DATAI_3_),
.Z(U3349));
MUX2_X1 U9385 (.S(U3149),
.A(n11369),
.B(DATAI_2_),
.Z(U3350));
MUX2_X1 U9386 (.S(U3149),
.A(n13778),
.B(DATAI_1_),
.Z(U3351));
OAI22_X1 U9387 (.B2(n13779),
.B1(n13780),
.A1(n13782),
.A2(n13781),
.ZN(n13783));
AOI21_X1 U9388 (.A(n13783),
.B2(n13784),
.B1(n13785),
.ZN(n13786));
OAI21_X1 U9389 (.A(n13786),
.B2(n13787),
.B1(n13844),
.ZN(n13788));
AOI21_X1 U9390 (.A(n13788),
.B2(n13789),
.B1(n13790),
.ZN(n13791));
OAI21_X1 U9391 (.A(n13791),
.B2(n13792),
.B1(n11157),
.ZN(U3286));
INV_X1 U9393 (.A(n13805),
.ZN(n13797));
INV_X1 U9394 (.A(n13794),
.ZN(n13800));
NOR3_X1 U9395 (.A3(n13795),
.A1(n13800),
.A2(n13799),
.ZN(n13796));
AOI21_X1 U9396 (.A(n13796),
.B2(n13804),
.B1(n13797),
.ZN(n13809));
OAI21_X1 U9397 (.A(n13798),
.B2(n13799),
.B1(n13800),
.ZN(n13802));
NAND2_X1 U9398 (.A2(n13801),
.A1(n13802),
.ZN(n13803));
AOI21_X1 U9399 (.A(n13803),
.B2(n13804),
.B1(n13805),
.ZN(n13808));
AOI22_X1 U9400 (.B2(U3149),
.B1(REG3_REG_17__SCAN_IN),
.A1(ADDR_REG_17__SCAN_IN),
.A2(FE_OFN1_n13320),
.ZN(n13807));
OAI221_X1 U9401 (.C2(n13808),
.C1(n13812),
.A(n13807),
.B2(n13809),
.B1(n13810),
.ZN(U3257));
INV_X1 U9402 (.A(DATAI_17_),
.ZN(n13811));
AOI22_X1 U9403 (.B2(U3149),
.B1(n13811),
.A1(STATE_REG_SCAN_IN),
.A2(n13812),
.ZN(U3335));
OAI22_X1 U9404 (.B2(STATE_REG_SCAN_IN),
.B1(DATAI_0_),
.A1(U3149),
.A2(IR_REG_0__SCAN_IN),
.ZN(n13813));
INV_X1 U9405 (.A(n13813),
.ZN(U3352));
AND2_X1 U9406 (.A2(n13814),
.A1(D_REG_31__SCAN_IN),
.ZN(U3291));
AND2_X1 U9407 (.A2(n13814),
.A1(D_REG_30__SCAN_IN),
.ZN(U3292));
AND2_X1 U9408 (.A2(n13814),
.A1(D_REG_29__SCAN_IN),
.ZN(U3293));
AND2_X1 U9409 (.A2(n13814),
.A1(D_REG_28__SCAN_IN),
.ZN(U3294));
AND2_X1 U9410 (.A2(n13814),
.A1(D_REG_27__SCAN_IN),
.ZN(U3295));
AND2_X1 U9411 (.A2(n13814),
.A1(D_REG_26__SCAN_IN),
.ZN(U3296));
AND2_X1 U9412 (.A2(n13814),
.A1(D_REG_25__SCAN_IN),
.ZN(U3297));
AND2_X1 U9413 (.A2(n13814),
.A1(D_REG_24__SCAN_IN),
.ZN(U3298));
AND2_X1 U9414 (.A2(n13814),
.A1(D_REG_23__SCAN_IN),
.ZN(U3299));
AND2_X1 U9415 (.A2(n13814),
.A1(D_REG_22__SCAN_IN),
.ZN(U3300));
AND2_X1 U9416 (.A2(n13814),
.A1(D_REG_21__SCAN_IN),
.ZN(U3301));
AND2_X1 U9417 (.A2(n13814),
.A1(D_REG_20__SCAN_IN),
.ZN(U3302));
AND2_X1 U9418 (.A2(n13814),
.A1(D_REG_19__SCAN_IN),
.ZN(U3303));
AND2_X1 U9419 (.A2(n13814),
.A1(D_REG_18__SCAN_IN),
.ZN(U3304));
AND2_X1 U9420 (.A2(n13814),
.A1(D_REG_17__SCAN_IN),
.ZN(U3305));
AND2_X1 U9421 (.A2(n13814),
.A1(D_REG_16__SCAN_IN),
.ZN(U3306));
AND2_X1 U9422 (.A2(n13814),
.A1(D_REG_15__SCAN_IN),
.ZN(U3307));
AND2_X1 U9423 (.A2(n13814),
.A1(D_REG_14__SCAN_IN),
.ZN(U3308));
AND2_X1 U9424 (.A2(n13814),
.A1(D_REG_13__SCAN_IN),
.ZN(U3309));
AND2_X1 U9425 (.A2(n13814),
.A1(D_REG_12__SCAN_IN),
.ZN(U3310));
AND2_X1 U9426 (.A2(n13814),
.A1(D_REG_11__SCAN_IN),
.ZN(U3311));
AND2_X1 U9427 (.A2(n13814),
.A1(D_REG_10__SCAN_IN),
.ZN(U3312));
AND2_X1 U9428 (.A2(n13814),
.A1(D_REG_9__SCAN_IN),
.ZN(U3313));
AND2_X1 U9429 (.A2(n13814),
.A1(D_REG_8__SCAN_IN),
.ZN(U3314));
AND2_X1 U9430 (.A2(n13814),
.A1(D_REG_7__SCAN_IN),
.ZN(U3315));
AND2_X1 U9431 (.A2(n13814),
.A1(D_REG_6__SCAN_IN),
.ZN(U3316));
AND2_X1 U9432 (.A2(n13814),
.A1(D_REG_5__SCAN_IN),
.ZN(U3317));
AND2_X1 U9433 (.A2(n13814),
.A1(D_REG_4__SCAN_IN),
.ZN(U3318));
AND2_X1 U9434 (.A2(n13814),
.A1(D_REG_3__SCAN_IN),
.ZN(U3319));
AND2_X1 U9435 (.A2(n13814),
.A1(D_REG_2__SCAN_IN),
.ZN(U3320));
INV_X1 U9436 (.A(DATAI_23_),
.ZN(n13816));
OAI21_X1 U9437 (.A(n13815),
.B2(n13816),
.B1(STATE_REG_SCAN_IN),
.ZN(U3329));
AOI22_X1 U9438 (.B2(n13860),
.B1(n11359),
.A1(FE_OFN3_n13832),
.A2(n13817),
.ZN(U3467));
NOR2_X1 U9439 (.A2(n13818),
.A1(n13819),
.ZN(n13821));
AOI211_X1 U9440 (.C1(n13822),
.A(n13821),
.C2(n13829),
.B(n13820),
.ZN(n13838));
OAI22_X1 U9441 (.B2(n13823),
.B1(FE_OFN3_n13832),
.A1(FE_OFN21_n13759),
.A2(n13834),
.ZN(n13825));
INV_X1 U9442 (.A(n13825),
.ZN(n13826));
OAI21_X1 U9443 (.A(n13826),
.B2(n13860),
.B1(n13838),
.ZN(U3477));
AOI211_X1 U9444 (.C1(n13830),
.A(n13828),
.C2(n13829),
.B(n13827),
.ZN(n13840));
AOI22_X1 U9445 (.B2(n13860),
.B1(n11405),
.A1(FE_OFN3_n13832),
.A2(n13840),
.ZN(U3479));
OAI22_X1 U9446 (.B2(n13833),
.B1(n13841),
.A1(FE_OFN7_n13835),
.A2(n13834),
.ZN(n13836));
INV_X1 U9447 (.A(n13836),
.ZN(n13837));
OAI21_X1 U9448 (.A(n13837),
.B2(n13839),
.B1(n13838),
.ZN(U3523));
AOI22_X1 U9449 (.B2(n13839),
.B1(n11409),
.A1(n13841),
.A2(n13840),
.ZN(U3524));
AOI22_X1 U9450 (.B2(n13842),
.B1(REG3_REG_2__SCAN_IN),
.A1(REG2_REG_2__SCAN_IN),
.A2(n11157),
.ZN(n13849));
OAI22_X1 U9451 (.B2(n13843),
.B1(n13844),
.A1(n13846),
.A2(n13845),
.ZN(n13847));
INV_X1 U9452 (.A(n13847),
.ZN(n13848));
OAI211_X1 U9453 (.C1(n11157),
.A(n13849),
.C2(n13850),
.B(n13848),
.ZN(U3288));
OAI21_X1 U6520 (.A(n13853),
.B2(n12155),
.B1(n13860),
.ZN(U3514));
INV_X1 U6530 (.A(n12016),
.ZN(n13853));
OAI211_X1 U6550 (.C1(n13839),
.A(n12152),
.C2(n12150),
.B(n11306),
.ZN(U3543));
OAI211_X1 U6556 (.C1(n12157),
.A(n12117),
.C2(n13844),
.B(n12121),
.ZN(U3262));
OAI21_X1 U6557 (.A(n13854),
.B2(n13115),
.B1(n11816),
.ZN(n11828));
AOI21_X1 U6564 (.A(n13584),
.B2(n13115),
.B1(n11816),
.ZN(n13854));
INV_X1 U6568 (.A(n13789),
.ZN(n13584));
INV_X1 U6570 (.A(n12204),
.ZN(n12214));
NAND2_X1 U6572 (.A2(n12198),
.A1(STATE_REG_SCAN_IN),
.ZN(n12204));
INV_X1 U6575 (.A(n13855),
.ZN(n12569));
OAI21_X1 U6600 (.A(n12633),
.B2(n12680),
.B1(n13779),
.ZN(n13855));
INV_X1 U6604 (.A(n13856),
.ZN(n12070));
OAI21_X1 U6605 (.A(n12067),
.B2(n13014),
.B1(n12132),
.ZN(n13856));
AOI211_X1 U6609 (.C1(n13016),
.A(n12081),
.C2(n13361),
.B(n13857),
.ZN(n12084));
NOR2_X1 U6617 (.A2(n13355),
.A1(n13014),
.ZN(n13857));
AOI21_X1 U6619 (.A(n13858),
.B2(n13839),
.B1(REG1_REG_27__SCAN_IN),
.ZN(n12148));
NOR2_X1 U6620 (.A2(n13325),
.A1(FE_OFN7_n13835),
.ZN(n13858));
AOI21_X1 U6622 (.A(n13859),
.B2(n13729),
.B1(n11803),
.ZN(n11308));
NOR2_X1 U6623 (.A2(FE_OFN3_n13832),
.A1(n11804),
.ZN(n13859));
INV_X4 U6629 (.A(n13223),
.ZN(U4043));
NAND2_X1 U6658 (.A2(n12167),
.A1(n12170),
.ZN(n13223));
NAND2_X2 U6675 (.A2(n13846),
.A1(n11819),
.ZN(n13789));
INV_X1 U6676 (.A(REG1_REG_6__SCAN_IN),
.ZN(n11409));
XNOR2_X1 U6681 (.B(n12320),
.A(REG1_REG_6__SCAN_IN),
.ZN(n12284));
OAI22_X1 U6683 (.B2(n12282),
.B1(n12283),
.A1(n13775),
.A2(REG1_REG_5__SCAN_IN),
.ZN(n12320));
XNOR2_X1 U6685 (.B(n12771),
.A(n12772),
.ZN(n12582));
OAI21_X1 U6690 (.A(n12581),
.B2(n11194),
.B1(n12661),
.ZN(n12771));
INV_X1 U6691 (.A(REG1_REG_15__SCAN_IN),
.ZN(n12772));
OR2_X1 U6692 (.A2(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN),
.A1(n12776),
.ZN(n12778));
OR2_X1 U6694 (.A2(n12935),
.A1(n13014),
.ZN(n12098));
AOI21_X1 U6695 (.A(n11648),
.B2(n11644),
.B1(n13328),
.ZN(n12935));
INV_X1 U6698 (.A(n13035),
.ZN(n13014));
INV_X1 U6701 (.A(n12237),
.ZN(n13078));
NAND2_X1 U6702 (.A2(n13124),
.A1(n13122),
.ZN(n12237));
INV_X1 U6705 (.A(n11271),
.ZN(n12040));
NAND2_X1 U6711 (.A2(n12129),
.A1(n11272),
.ZN(n11271));
INV_X1 U6712 (.A(n13860),
.ZN(n13832));
NAND2_X2 U6725 (.A2(n12027),
.A1(n13918),
.ZN(n13860));
NAND2_X1 U6726 (.A2(n13860),
.A1(REG0_REG_28__SCAN_IN),
.ZN(n12015));
XNOR2_X1 U6731 (.B(n12379),
.A(n12642),
.ZN(n12374));
NAND2_X1 U6733 (.A2(n11431),
.A1(n11446),
.ZN(n12379));
INV_X1 U6734 (.A(REG1_REG_7__SCAN_IN),
.ZN(n12642));
XNOR2_X1 U6736 (.B(n13288),
.A(n13275),
.ZN(n12770));
NAND2_X1 U6738 (.A2(n11514),
.A1(n11567),
.ZN(n13288));
INV_X1 U6745 (.A(REG2_REG_16__SCAN_IN),
.ZN(n13275));
XNOR2_X1 U6747 (.B(n12240),
.A(n12498),
.ZN(n12186));
NAND2_X1 U6749 (.A2(n12178),
.A1(n13227),
.ZN(n12240));
INV_X1 U6753 (.A(REG2_REG_3__SCAN_IN),
.ZN(n12498));
XNOR2_X1 U6767 (.B(n13793),
.A(n13653),
.ZN(n13805));
NAND2_X1 U6769 (.A2(n13290),
.A1(n13289),
.ZN(n13793));
INV_X1 U6774 (.A(REG1_REG_17__SCAN_IN),
.ZN(n13653));
INV_X1 U6775 (.A(n12848),
.ZN(n13196));
NAND2_X1 U6782 (.A2(n11569),
.A1(DATAI_30_),
.ZN(n12848));
INV_X1 U6785 (.A(n12903),
.ZN(n13537));
NAND2_X1 U6787 (.A2(n11526),
.A1(n11525),
.ZN(n12903));
INV_X1 U6788 (.A(n12091),
.ZN(n13861));
NOR2_X1 U6789 (.A2(n13861),
.A1(n12090),
.ZN(n11310));
INV_X1 U6790 (.A(n12060),
.ZN(n13862));
NOR2_X1 U6791 (.A2(n13862),
.A1(n12059),
.ZN(n11311));
INV_X1 U6805 (.A(n12075),
.ZN(n13863));
NOR2_X1 U6815 (.A2(n13863),
.A1(n12074),
.ZN(n11303));
INV_X1 U6821 (.A(n12104),
.ZN(n13864));
NOR2_X1 U6829 (.A2(n13864),
.A1(n12103),
.ZN(n11312));
XNOR2_X1 U6835 (.B(n13430),
.A(n13869),
.ZN(n13637));
NAND2_X1 U6839 (.A2(n13421),
.A1(n13420),
.ZN(n13430));
INV_X1 U6840 (.A(n13865),
.ZN(n12157));
AOI21_X1 U6842 (.A(n12012),
.B2(n12051),
.B1(n12932),
.ZN(n13865));
INV_X1 U6845 (.A(n11800),
.ZN(n12012));
AOI21_X1 U6846 (.A(n13533),
.B2(n13531),
.B1(n13530),
.ZN(n13676));
NOR2_X1 U6847 (.A2(n13530),
.A1(n13531),
.ZN(n13533));
INV_X2 U6848 (.A(n13795),
.ZN(n13798));
NAND2_X2 U6850 (.A2(n12227),
.A1(n12174),
.ZN(n13795));
INV_X2 U6852 (.A(n13016),
.ZN(n13041));
NAND2_X1 U6859 (.A2(n11992),
.A1(n13815),
.ZN(n13016));
OAI211_X1 U6861 (.C1(n13404),
.A(n13672),
.C2(n13417),
.B(n13866),
.ZN(n13626));
NAND2_X1 U6864 (.A2(n13417),
.A1(n13404),
.ZN(n13866));
NAND2_X2 U6867 (.A2(n11685),
.A1(n13193),
.ZN(n13672));
OR2_X1 U6871 (.A2(n13633),
.A1(n13431),
.ZN(n13432));
XOR2_X1 U6873 (.B(n12444),
.A(n13083),
.Z(n12451));
NAND2_X1 U6876 (.A2(n11697),
.A1(n11696),
.ZN(n12444));
INV_X1 U6890 (.A(n12813),
.ZN(n13867));
NOR2_X1 U6891 (.A2(n13867),
.A1(n12812),
.ZN(n12815));
NOR2_X1 U6904 (.A2(n11812),
.A1(n13919),
.ZN(n13580));
AOI21_X1 U6907 (.A(n12438),
.B2(n12439),
.B1(n12490),
.ZN(n12496));
NOR2_X1 U6908 (.A2(n12490),
.A1(n12439),
.ZN(n12438));
AOI21_X1 U6909 (.A(n11282),
.B2(n11279),
.B1(n11175),
.ZN(n13869));
OAI21_X1 U6912 (.A(n13870),
.B2(n12556),
.B1(n13099),
.ZN(n12633));
AOI21_X1 U6915 (.A(n13568),
.B2(n12556),
.B1(n13099),
.ZN(n13870));
INV_X2 U6916 (.A(n13577),
.ZN(n13785));
NAND2_X1 U6919 (.A2(n13782),
.A1(n13688),
.ZN(n13577));
INV_X2 U6923 (.A(n13292),
.ZN(n13801));
NOR2_X2 U6924 (.A2(n12182),
.A1(n13764),
.ZN(n13292));
XNOR2_X1 U6926 (.B(n12571),
.A(n13704),
.ZN(n12403));
OAI21_X1 U6927 (.A(n12395),
.B2(n11191),
.B1(n13239),
.ZN(n12571));
INV_X1 U6928 (.A(REG1_REG_11__SCAN_IN),
.ZN(n13704));
INV_X1 U6930 (.A(n13598),
.ZN(n13871));
AOI21_X1 U6931 (.A(n13596),
.B2(n13829),
.B1(n13871),
.ZN(n13600));
XOR2_X1 U6932 (.B(n12561),
.A(n13099),
.Z(n12631));
NAND2_X1 U6933 (.A2(n11710),
.A1(n11709),
.ZN(n12561));
XOR2_X1 U6936 (.B(n13872),
.A(n13448),
.Z(n13645));
NAND2_X1 U6939 (.A2(n11280),
.A1(n11728),
.ZN(n13872));
NAND2_X1 U6940 (.A2(n12944),
.A1(n11248),
.ZN(n11247));
OR2_X1 U6949 (.A2(n11954),
.A1(n11953),
.ZN(n12944));
NAND2_X1 U6951 (.A2(n11945),
.A1(n12982),
.ZN(n11248));
NAND2_X1 U6952 (.A2(n12011),
.A1(n11799),
.ZN(n11800));
INV_X1 U6964 (.A(n11245),
.ZN(n12234));
NAND2_X1 U6974 (.A2(n13091),
.A1(n11838),
.ZN(n11245));
OAI21_X1 U6975 (.A(n13424),
.B2(n13422),
.B1(n13423),
.ZN(n13446));
NAND2_X1 U6976 (.A2(n11915),
.A1(n12976),
.ZN(n13424));
INV_X1 U6985 (.A(n13873),
.ZN(n12045));
AOI22_X1 U6986 (.B2(n13210),
.B1(n13690),
.A1(n13688),
.A2(n13212),
.ZN(n13873));
AOI22_X1 U6987 (.B2(n13874),
.B1(n13876),
.A1(n13307),
.A2(n13879),
.ZN(n13305));
OR2_X1 U6989 (.A2(n13879),
.A1(n13307),
.ZN(n13874));
INV_X1 U7000 (.A(n11687),
.ZN(n13875));
NAND2_X1 U7002 (.A2(B_REG_SCAN_IN),
.A1(n13875),
.ZN(n11689));
OAI21_X1 U7007 (.A(n13368),
.B2(n11737),
.B1(n11736),
.ZN(n13598));
NAND2_X1 U7008 (.A2(n11737),
.A1(n11736),
.ZN(n13368));
INV_X1 U7010 (.A(n13302),
.ZN(n13876));
OAI22_X1 U7012 (.B2(n13291),
.B1(n13793),
.A1(n13653),
.A2(n13812),
.ZN(n13302));
INV_X1 U7036 (.A(n11248),
.ZN(n12984));
NAND2_X1 U7060 (.A2(n13877),
.A1(n13059),
.ZN(n11210));
INV_X1 U7083 (.A(n12042),
.ZN(n13877));
NAND2_X1 U7084 (.A2(n11641),
.A1(n13060),
.ZN(n12042));
INV_X1 U7104 (.A(n11944),
.ZN(n12943));
NOR2_X1 U7105 (.A2(n12982),
.A1(n11945),
.ZN(n11944));
INV_X1 U7112 (.A(n13878),
.ZN(n13379));
AOI21_X1 U7114 (.A(n13376),
.B2(n13377),
.B1(n13375),
.ZN(n13878));
INV_X2 U7115 (.A(n13819),
.ZN(n13688));
NAND2_X2 U7116 (.A2(n12168),
.A1(n13764),
.ZN(n13819));
INV_X1 U7124 (.A(REG1_REG_18__SCAN_IN),
.ZN(n13879));
NAND2_X1 U7125 (.A2(n11556),
.A1(n12212),
.ZN(n13307));
NOR3_X1 U7127 (.A3(n12172),
.A1(n12189),
.A2(n13880),
.ZN(n12227));
INV_X1 U7137 (.A(n12190),
.ZN(n13880));
NAND2_X1 U7138 (.A2(n12168),
.A1(n12170),
.ZN(n12190));
NAND3_X1 U7139 (.A3(n11808),
.A1(n13881),
.A2(n11990),
.ZN(n12028));
INV_X1 U7142 (.A(n11812),
.ZN(n13881));
NAND2_X1 U7144 (.A2(n13203),
.A1(n11789),
.ZN(n11812));
INV_X1 U7145 (.A(n11273),
.ZN(n12125));
NOR2_X1 U7150 (.A2(n13343),
.A1(n12889),
.ZN(n11273));
INV_X1 U7151 (.A(n13184),
.ZN(n13180));
NAND2_X1 U7152 (.A2(n13059),
.A1(n13060),
.ZN(n13184));
INV_X1 U7153 (.A(n13882),
.ZN(n12908));
AOI22_X1 U7154 (.B2(n13640),
.B1(n11846),
.A1(FE_OFN0_n11847),
.A2(n13438),
.ZN(n13882));
INV_X1 U7156 (.A(n12453),
.ZN(n13662));
NAND3_X1 U7157 (.A3(n11838),
.A1(n13769),
.A2(n13189),
.ZN(n12453));
AOI211_X1 U7160 (.C1(n13279),
.A(n13280),
.C2(n13278),
.B(REG2_REG_17__SCAN_IN),
.ZN(n13799));
INV_X1 U7162 (.A(n11945),
.ZN(n12988));
NAND2_X1 U7164 (.A2(n11942),
.A1(n11941),
.ZN(n11945));
INV_X1 U7166 (.A(n13066),
.ZN(n13065));
NOR2_X1 U7168 (.A2(n13209),
.A1(n11801),
.ZN(n13066));
INV_X1 U7172 (.A(n13375),
.ZN(n13350));
NAND2_X1 U7173 (.A2(n13628),
.A1(n13611),
.ZN(n13375));
OAI211_X1 U7185 (.C1(n13280),
.A(n13278),
.C2(n13279),
.B(REG2_REG_17__SCAN_IN),
.ZN(n13794));
INV_X1 U7187 (.A(n12314),
.ZN(n13204));
NAND3_X1 U7192 (.A3(STATE_REG_SCAN_IN),
.A1(n12166),
.A2(n12170),
.ZN(n12314));
INV_X1 U7193 (.A(n12126),
.ZN(n12124));
NAND2_X1 U7194 (.A2(n13343),
.A1(n12889),
.ZN(n12126));
INV_X1 U7219 (.A(n13324),
.ZN(n11974));
NAND2_X1 U7231 (.A2(n11569),
.A1(DATAI_27_),
.ZN(n13324));
OAI21_X1 U7236 (.A(n13883),
.B2(n11825),
.B1(FE_OFN16_n11466),
.ZN(n13209));
INV_X1 U7249 (.A(n11667),
.ZN(n13883));
OAI21_X1 U7271 (.A(n13884),
.B2(n11786),
.B1(n11787),
.ZN(n11984));
INV_X1 U7273 (.A(n12222),
.ZN(n13884));
NAND2_X1 U7287 (.A2(n11767),
.A1(n13766),
.ZN(n12222));
INV_X1 U7292 (.A(n13085),
.ZN(n13423));
NAND2_X1 U7299 (.A2(n13656),
.A1(n13471),
.ZN(n13085));
INV_X1 U7301 (.A(n13092),
.ZN(n13090));
AOI22_X1 U7302 (.B2(n13196),
.B1(n13197),
.A1(n13208),
.A2(n13069),
.ZN(n13092));
NAND2_X1 U7315 (.A2(n11776),
.A1(n11775),
.ZN(n12170));
OAI21_X1 U7328 (.A(n12771),
.B2(n12773),
.B1(n12772),
.ZN(n12775));
INV_X1 U7329 (.A(n12032),
.ZN(n12877));
NAND2_X1 U7330 (.A2(n11569),
.A1(DATAI_26_),
.ZN(n12032));
INV_X1 U7331 (.A(n11736),
.ZN(n13366));
NAND2_X1 U7332 (.A2(n13121),
.A1(n13175),
.ZN(n11736));
AOI21_X1 U7348 (.A(n13885),
.B2(n12141),
.B1(n13343),
.ZN(n12019));
INV_X1 U7349 (.A(n13072),
.ZN(n13885));
NAND2_X1 U7351 (.A2(n13213),
.A1(n13337),
.ZN(n13072));
OAI21_X2 U7364 (.A(n13886),
.B2(n12880),
.B1(FE_OFN16_n11466),
.ZN(n13212));
INV_X1 U7387 (.A(n11627),
.ZN(n13886));
INV_X1 U7426 (.A(n13395),
.ZN(n13611));
NAND2_X1 U7428 (.A2(n11569),
.A1(DATAI_21_),
.ZN(n13395));
INV_X1 U7431 (.A(n13427),
.ZN(n13612));
AOI21_X1 U7432 (.A(n11577),
.B2(n11644),
.B1(n13409),
.ZN(n13427));
AOI21_X1 U7439 (.A(n13889),
.B2(n11994),
.B1(n11642),
.ZN(n13328));
INV_X1 U7445 (.A(n13889),
.ZN(n11654));
NOR2_X1 U7474 (.A2(n11642),
.A1(n11994),
.ZN(n13889));
OAI21_X1 U7482 (.A(n12662),
.B2(n13770),
.B1(REG2_REG_14__SCAN_IN),
.ZN(n12593));
OAI22_X1 U7486 (.B2(n12590),
.B1(n13264),
.A1(n13269),
.A2(n12589),
.ZN(n12662));
INV_X1 U7491 (.A(n13213),
.ZN(n13355));
NAND2_X1 U7493 (.A2(n11620),
.A1(n11619),
.ZN(n13213));
INV_X1 U7494 (.A(n13890),
.ZN(n13343));
AOI21_X1 U7495 (.A(n11636),
.B2(n12064),
.B1(n11644),
.ZN(n13890));
OAI21_X2 U7496 (.A(n13891),
.B2(n13398),
.B1(FE_OFN16_n11466),
.ZN(n13605));
INV_X1 U7502 (.A(n11605),
.ZN(n13891));
AOI21_X2 U7507 (.A(n11596),
.B2(n13381),
.B1(n11644),
.ZN(n13614));
NAND2_X1 U7518 (.A2(n13920),
.A1(n13482),
.ZN(n13164));
AOI21_X1 U7537 (.A(n13894),
.B2(n13445),
.B1(n13420),
.ZN(n11572));
INV_X1 U7566 (.A(n13894),
.ZN(n13421));
NOR2_X1 U7572 (.A2(n13640),
.A1(n13633),
.ZN(n13894));
INV_X1 U7574 (.A(n11728),
.ZN(n13895));
NOR2_X1 U7575 (.A2(n13895),
.A1(n11730),
.ZN(n11175));
NOR2_X1 U7576 (.A2(n13896),
.A1(n11587),
.ZN(n13341));
NOR2_X1 U7578 (.A2(n12079),
.A1(FE_OFN16_n11466),
.ZN(n13896));
OAI21_X1 U7581 (.A(n12584),
.B2(n13771),
.B1(REG2_REG_11__SCAN_IN),
.ZN(n12586));
OAI21_X1 U7586 (.A(n13900),
.B2(n13240),
.B1(n12400),
.ZN(n12584));
INV_X1 U7587 (.A(n13897),
.ZN(n11436));
OAI21_X1 U7605 (.A(n13087),
.B2(n13899),
.B1(n12526),
.ZN(n13897));
OAI21_X2 U7612 (.A(n13898),
.B2(n13473),
.B1(FE_OFN16_n11466),
.ZN(n13656));
INV_X1 U7613 (.A(n11564),
.ZN(n13898));
INV_X1 U7616 (.A(n13139),
.ZN(n13899));
NAND2_X1 U7617 (.A2(n13772),
.A1(REG2_REG_10__SCAN_IN),
.ZN(n13900));
INV_X1 U7629 (.A(n13689),
.ZN(n13525));
NAND4_X1 U7644 (.A4(n11501),
.A3(n11504),
.A1(n11503),
.A2(n11502),
.ZN(n13689));
INV_X1 U7677 (.A(n11294),
.ZN(n11296));
NAND2_X1 U7697 (.A2(n11863),
.A1(n12629),
.ZN(n11294));
INV_X1 U7714 (.A(n13217),
.ZN(n12828));
NAND4_X1 U7715 (.A4(n11442),
.A3(n11443),
.A1(n11444),
.A2(n11445),
.ZN(n13217));
INV_X1 U7716 (.A(n13655),
.ZN(n13526));
NAND3_X1 U7723 (.A3(n11522),
.A1(n11521),
.A2(n11520),
.ZN(n13655));
INV_X1 U7725 (.A(n13666),
.ZN(n13545));
NAND4_X1 U7726 (.A4(n11529),
.A3(n11528),
.A1(n11531),
.A2(n11530),
.ZN(n13666));
INV_X1 U7729 (.A(n13219),
.ZN(n12652));
NAND4_X1 U7740 (.A4(n11413),
.A3(n11412),
.A1(n11410),
.A2(n11411),
.ZN(n13219));
INV_X1 U7743 (.A(n13218),
.ZN(n12675));
NAND4_X1 U7748 (.A4(n11423),
.A3(n11426),
.A1(n11425),
.A2(n11424),
.ZN(n13218));
AOI21_X1 U7751 (.A(n13901),
.B2(n11498),
.B1(n11499),
.ZN(n13551));
INV_X1 U7758 (.A(n13901),
.ZN(n11187));
NOR2_X1 U7760 (.A2(n11499),
.A1(n11498),
.ZN(n13901));
NAND2_X1 U7853 (.A2(REG2_REG_14__SCAN_IN),
.A1(FE_OFN27_n11469),
.ZN(n11529));
INV_X1 U7907 (.A(n13903),
.ZN(n12349));
AOI211_X1 U7908 (.C1(n12372),
.A(n12325),
.C2(n12324),
.B(REG1_REG_8__SCAN_IN),
.ZN(n13903));
INV_X1 U7909 (.A(n13904),
.ZN(n12356));
AOI22_X1 U7915 (.B2(n12377),
.B1(n12333),
.A1(REG2_REG_7__SCAN_IN),
.A2(n12334),
.ZN(n13904));
OAI21_X1 U7918 (.A(n13905),
.B2(n12320),
.B1(n11409),
.ZN(n12372));
NAND2_X1 U7919 (.A2(n12319),
.A1(n13774),
.ZN(n13905));
INV_X1 U7921 (.A(WxUoeaFQeyYVaGStCqAbTWICyXpTFvtD_Z),
.ZN(n12357));
NAND2_X1 U7926 (.A2(n11449),
.A1(n11495),
.ZN(n12354));
NAND2_X1 U7991 (.A2(REG2_REG_9__SCAN_IN),
.A1(FE_DBTN0_n11469),
.ZN(n11460));
OAI21_X1 U7993 (.A(n11464),
.B2(n11207),
.B1(REG3_REG_9__SCAN_IN),
.ZN(n12760));
NAND2_X1 U7994 (.A2(n11207),
.A1(REG3_REG_9__SCAN_IN),
.ZN(n11464));
INV_X1 U7995 (.A(n13907),
.ZN(n11791));
AOI22_X1 U8028 (.B2(n12196),
.B1(n11761),
.A1(IR_REG_24__SCAN_IN),
.A2(n12198),
.ZN(n12138));
INV_X1 U8035 (.A(n13908),
.ZN(n12377));
AOI22_X1 U8040 (.B2(n12330),
.B1(n12329),
.A1(REG2_REG_6__SCAN_IN),
.A2(n13774),
.ZN(n13908));
NAND2_X1 U8047 (.A2(REG2_REG_10__SCAN_IN),
.A1(FE_DBTN0_n11469),
.ZN(n11470));
NAND2_X1 U8059 (.A2(REG2_REG_2__SCAN_IN),
.A1(FE_DBTN0_n11469),
.ZN(n11373));
OAI21_X1 U8073 (.A(IR_REG_21__SCAN_IN),
.B2(n11676),
.B1(n12198),
.ZN(n11680));
NAND2_X1 U8076 (.A2(FE_DBTN1_n11467),
.A1(REG1_REG_1__SCAN_IN),
.ZN(n11346));
NAND2_X1 U8078 (.A2(n11341),
.A1(n13763),
.ZN(n11467));
NAND2_X1 U8089 (.A2(REG2_REG_1__SCAN_IN),
.A1(FE_DBTN0_n11469),
.ZN(n11345));
NAND3_X1 U8095 (.A3(REG3_REG_9__SCAN_IN),
.A1(n11207),
.A2(REG3_REG_10__SCAN_IN),
.ZN(n11475));
NOR2_X1 U8096 (.A2(n11439),
.A1(n11438),
.ZN(n11207));
INV_X1 U8099 (.A(n13913),
.ZN(n11363));
OAI22_X1 U8105 (.B2(n11418),
.B1(n11359),
.A1(n12551),
.A2(n11469),
.ZN(n13913));
INV_X1 U8106 (.A(n11207),
.ZN(n11454));
NAND3_X1 U8107 (.A3(n13914),
.A1(n12243),
.A2(n13781),
.ZN(n12272));
NAND2_X1 U8114 (.A2(n12242),
.A1(n12241),
.ZN(n13914));
AOI211_X1 U8120 (.C1(IR_REG_31__SCAN_IN),
.A(n13916),
.C2(IR_REG_27__SCAN_IN),
.B(n13915),
.ZN(n11288));
INV_X1 U8122 (.A(n11289),
.ZN(n13915));
AOI21_X1 U8136 (.A(n13917),
.B2(IR_REG_26__SCAN_IN),
.B1(IR_REG_31__SCAN_IN),
.ZN(n11289));
INV_X1 U8139 (.A(n11391),
.ZN(n11389));
NOR2_X1 U8181 (.A2(n11171),
.A1(IR_REG_3__SCAN_IN),
.ZN(n11391));
OR2_X1 U8182 (.A2(REG1_REG_2__SCAN_IN),
.A1(n12179),
.ZN(n13225));
INV_X1 U8196 (.A(n12248),
.ZN(n13776));
NAND2_X1 U8197 (.A2(n11380),
.A1(n11389),
.ZN(n12248));
INV_X1 U8198 (.A(IR_REG_28__SCAN_IN),
.ZN(n13916));
INV_X1 U8228 (.A(n11347),
.ZN(n13917));
OR2_X1 U8261 (.A2(REG2_REG_2__SCAN_IN),
.A1(n12175),
.ZN(n13227));
INV_X1 U8262 (.A(IR_REG_25__SCAN_IN),
.ZN(n11329));
NOR3_X1 U8266 (.A3(IR_REG_25__SCAN_IN),
.A1(n11330),
.A2(IR_REG_29__SCAN_IN),
.ZN(n11258));
INV_X1 U8267 (.A(n12028),
.ZN(n13918));
NAND2_X1 U6526 (.A2(n13153),
.A1(n13154),
.ZN(n11186));
AOI21_X1 U6549 (.A(n11744),
.B2(n11745),
.B1(n11746),
.ZN(n12002));
NOR2_X1 U6632 (.A2(n11770),
.A1(n13907),
.ZN(n11772));
MUX2_X1 U6732 (.S(IR_REG_29__SCAN_IN),
.A(IR_REG_31__SCAN_IN),
.B(n11335),
.Z(n11337));
AND4_X1 U6903 (.A4(n11477),
.A3(n11478),
.A1(n11480),
.A2(n11479),
.ZN(n13578));
OR2_X1 U7388 (.A2(n11811),
.A1(n11983),
.ZN(n13919));
AND2_X1 U7411 (.A2(n13167),
.A1(n13485),
.ZN(n13920));
OR2_X1 U7440 (.A2(n12784),
.A1(n12785),
.ZN(n13921));
NAND4_X2 NreNGPwwSfGxuZEJRmMXTmzYADEemtnb (.A4(n13008),
.A3(n11689),
.A2(n13306),
.A1(n12395),
.ZN(NreNGPwwSfGxuZEJRmMXTmzYADEemtnb_ZN));
OR3_X1 qQydNHNCopcDTmEyGIIdyrFQIErIFgJX (.A3(n13090),
.A2(n13839),
.A1(n13565),
.ZN(qQydNHNCopcDTmEyGIIdyrFQIErIFgJX_ZN));
AOI22_X4 lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL (.B2(n12515),
.B1(n13129),
.A1(n13313),
.A2(n11495),
.ZN(lkXvcZHjgjWzZgjbcIpFrxTZHAjqZjhL_ZN));
OR2_X1 FzxTCFmmmorPYWBoKVOYVzYHHyJMkxJR (.A2(n12515),
.A1(n13491),
.ZN(FzxTCFmmmorPYWBoKVOYVzYHHyJMkxJR_ZN));
BUF_X1 rlUqTqnDczmjZLOdxrCVPPbsubqicwLv (.A(n13396),
.Z(rlUqTqnDczmjZLOdxrCVPPbsubqicwLv_Z));
NAND4_X2 KgXiNKYImGwoITNkFdnqdBmiQCHYgIoS (.A3(n11720),
.A4(n11824),
.A2(n12812),
.A1(n13611),
.ZN(KgXiNKYImGwoITNkFdnqdBmiQCHYgIoS_ZN));
BUF_X32 jexoRSiRmgnTTbxiBcsGLhbKTivhVojg (.A(n12362),
.Z(jexoRSiRmgnTTbxiBcsGLhbKTivhVojg_Z));
CLKBUF_X1 WxUoeaFQeyYVaGStCqAbTWICyXpTFvtD (.A(n12354),
.Z(WxUoeaFQeyYVaGStCqAbTWICyXpTFvtD_Z));

endmodule
